//Copyright (C)2014-2022 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//GOWIN Version: V1.9.8.07 Education
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9C
//Created Time: Wed Jan 04 22:52:53 2023

module Gowin_RAM16SDP (dout, wre, wad, di, rad, clk);

output [7:0] dout;
input wre;
input [9:0] wad;
input [7:0] di;
input [9:0] rad;
input clk;

wire wad4_inv;
wire wad5_inv;
wire wad6_inv;
wire lut_f_0;
wire wad7_inv;
wire wad8_inv;
wire wad9_inv;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire lut_f_20;
wire lut_f_21;
wire lut_f_22;
wire lut_f_23;
wire lut_f_24;
wire lut_f_25;
wire lut_f_26;
wire lut_f_27;
wire lut_f_28;
wire lut_f_29;
wire lut_f_30;
wire lut_f_31;
wire lut_f_32;
wire lut_f_33;
wire lut_f_34;
wire lut_f_35;
wire lut_f_36;
wire lut_f_37;
wire lut_f_38;
wire lut_f_39;
wire lut_f_40;
wire lut_f_41;
wire lut_f_42;
wire lut_f_43;
wire lut_f_44;
wire lut_f_45;
wire lut_f_46;
wire lut_f_47;
wire lut_f_48;
wire lut_f_49;
wire lut_f_50;
wire lut_f_51;
wire lut_f_52;
wire lut_f_53;
wire lut_f_54;
wire lut_f_55;
wire lut_f_56;
wire lut_f_57;
wire lut_f_58;
wire lut_f_59;
wire lut_f_60;
wire lut_f_61;
wire lut_f_62;
wire lut_f_63;
wire lut_f_64;
wire lut_f_65;
wire lut_f_66;
wire lut_f_67;
wire lut_f_68;
wire lut_f_69;
wire lut_f_70;
wire lut_f_71;
wire lut_f_72;
wire lut_f_73;
wire lut_f_74;
wire lut_f_75;
wire lut_f_76;
wire lut_f_77;
wire lut_f_78;
wire lut_f_79;
wire lut_f_80;
wire lut_f_81;
wire lut_f_82;
wire lut_f_83;
wire lut_f_84;
wire lut_f_85;
wire lut_f_86;
wire lut_f_87;
wire lut_f_88;
wire lut_f_89;
wire lut_f_90;
wire lut_f_91;
wire lut_f_92;
wire lut_f_93;
wire lut_f_94;
wire lut_f_95;
wire lut_f_96;
wire lut_f_97;
wire lut_f_98;
wire lut_f_99;
wire [3:0] ram16sdp_inst_0_dout;
wire [7:4] ram16sdp_inst_1_dout;
wire [3:0] ram16sdp_inst_2_dout;
wire [7:4] ram16sdp_inst_3_dout;
wire [3:0] ram16sdp_inst_4_dout;
wire [7:4] ram16sdp_inst_5_dout;
wire [3:0] ram16sdp_inst_6_dout;
wire [7:4] ram16sdp_inst_7_dout;
wire [3:0] ram16sdp_inst_8_dout;
wire [7:4] ram16sdp_inst_9_dout;
wire [3:0] ram16sdp_inst_10_dout;
wire [7:4] ram16sdp_inst_11_dout;
wire [3:0] ram16sdp_inst_12_dout;
wire [7:4] ram16sdp_inst_13_dout;
wire [3:0] ram16sdp_inst_14_dout;
wire [7:4] ram16sdp_inst_15_dout;
wire [3:0] ram16sdp_inst_16_dout;
wire [7:4] ram16sdp_inst_17_dout;
wire [3:0] ram16sdp_inst_18_dout;
wire [7:4] ram16sdp_inst_19_dout;
wire [3:0] ram16sdp_inst_20_dout;
wire [7:4] ram16sdp_inst_21_dout;
wire [3:0] ram16sdp_inst_22_dout;
wire [7:4] ram16sdp_inst_23_dout;
wire [3:0] ram16sdp_inst_24_dout;
wire [7:4] ram16sdp_inst_25_dout;
wire [3:0] ram16sdp_inst_26_dout;
wire [7:4] ram16sdp_inst_27_dout;
wire [3:0] ram16sdp_inst_28_dout;
wire [7:4] ram16sdp_inst_29_dout;
wire [3:0] ram16sdp_inst_30_dout;
wire [7:4] ram16sdp_inst_31_dout;
wire [3:0] ram16sdp_inst_32_dout;
wire [7:4] ram16sdp_inst_33_dout;
wire [3:0] ram16sdp_inst_34_dout;
wire [7:4] ram16sdp_inst_35_dout;
wire [3:0] ram16sdp_inst_36_dout;
wire [7:4] ram16sdp_inst_37_dout;
wire [3:0] ram16sdp_inst_38_dout;
wire [7:4] ram16sdp_inst_39_dout;
wire [3:0] ram16sdp_inst_40_dout;
wire [7:4] ram16sdp_inst_41_dout;
wire [3:0] ram16sdp_inst_42_dout;
wire [7:4] ram16sdp_inst_43_dout;
wire [3:0] ram16sdp_inst_44_dout;
wire [7:4] ram16sdp_inst_45_dout;
wire [3:0] ram16sdp_inst_46_dout;
wire [7:4] ram16sdp_inst_47_dout;
wire [3:0] ram16sdp_inst_48_dout;
wire [7:4] ram16sdp_inst_49_dout;
wire [3:0] ram16sdp_inst_50_dout;
wire [7:4] ram16sdp_inst_51_dout;
wire [3:0] ram16sdp_inst_52_dout;
wire [7:4] ram16sdp_inst_53_dout;
wire [3:0] ram16sdp_inst_54_dout;
wire [7:4] ram16sdp_inst_55_dout;
wire [3:0] ram16sdp_inst_56_dout;
wire [7:4] ram16sdp_inst_57_dout;
wire [3:0] ram16sdp_inst_58_dout;
wire [7:4] ram16sdp_inst_59_dout;
wire [3:0] ram16sdp_inst_60_dout;
wire [7:4] ram16sdp_inst_61_dout;
wire [3:0] ram16sdp_inst_62_dout;
wire [7:4] ram16sdp_inst_63_dout;
wire [3:0] ram16sdp_inst_64_dout;
wire [7:4] ram16sdp_inst_65_dout;
wire [3:0] ram16sdp_inst_66_dout;
wire [7:4] ram16sdp_inst_67_dout;
wire [3:0] ram16sdp_inst_68_dout;
wire [7:4] ram16sdp_inst_69_dout;
wire [3:0] ram16sdp_inst_70_dout;
wire [7:4] ram16sdp_inst_71_dout;
wire [3:0] ram16sdp_inst_72_dout;
wire [7:4] ram16sdp_inst_73_dout;
wire [3:0] ram16sdp_inst_74_dout;
wire [7:4] ram16sdp_inst_75_dout;
wire [3:0] ram16sdp_inst_76_dout;
wire [7:4] ram16sdp_inst_77_dout;
wire [3:0] ram16sdp_inst_78_dout;
wire [7:4] ram16sdp_inst_79_dout;
wire [3:0] ram16sdp_inst_80_dout;
wire [7:4] ram16sdp_inst_81_dout;
wire [3:0] ram16sdp_inst_82_dout;
wire [7:4] ram16sdp_inst_83_dout;
wire [3:0] ram16sdp_inst_84_dout;
wire [7:4] ram16sdp_inst_85_dout;
wire [3:0] ram16sdp_inst_86_dout;
wire [7:4] ram16sdp_inst_87_dout;
wire [3:0] ram16sdp_inst_88_dout;
wire [7:4] ram16sdp_inst_89_dout;
wire [3:0] ram16sdp_inst_90_dout;
wire [7:4] ram16sdp_inst_91_dout;
wire [3:0] ram16sdp_inst_92_dout;
wire [7:4] ram16sdp_inst_93_dout;
wire [3:0] ram16sdp_inst_94_dout;
wire [7:4] ram16sdp_inst_95_dout;
wire [3:0] ram16sdp_inst_96_dout;
wire [7:4] ram16sdp_inst_97_dout;
wire [3:0] ram16sdp_inst_98_dout;
wire [7:4] ram16sdp_inst_99_dout;
wire mux_o_0;
wire mux_o_1;
wire mux_o_2;
wire mux_o_3;
wire mux_o_4;
wire mux_o_5;
wire mux_o_6;
wire mux_o_7;
wire mux_o_8;
wire mux_o_9;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_17;
wire mux_o_18;
wire mux_o_19;
wire mux_o_20;
wire mux_o_21;
wire mux_o_22;
wire mux_o_23;
wire mux_o_24;
wire mux_o_25;
wire mux_o_26;
wire mux_o_27;
wire mux_o_28;
wire mux_o_29;
wire mux_o_30;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_38;
wire mux_o_39;
wire mux_o_40;
wire mux_o_41;
wire mux_o_42;
wire mux_o_43;
wire mux_o_45;
wire mux_o_46;
wire mux_o_47;
wire mux_o_49;
wire mux_o_50;
wire mux_o_52;
wire mux_o_53;
wire mux_o_54;
wire mux_o_55;
wire mux_o_56;
wire mux_o_57;
wire mux_o_58;
wire mux_o_59;
wire mux_o_60;
wire mux_o_61;
wire mux_o_62;
wire mux_o_63;
wire mux_o_64;
wire mux_o_65;
wire mux_o_66;
wire mux_o_67;
wire mux_o_68;
wire mux_o_69;
wire mux_o_70;
wire mux_o_71;
wire mux_o_72;
wire mux_o_73;
wire mux_o_74;
wire mux_o_75;
wire mux_o_76;
wire mux_o_77;
wire mux_o_78;
wire mux_o_79;
wire mux_o_80;
wire mux_o_81;
wire mux_o_82;
wire mux_o_83;
wire mux_o_84;
wire mux_o_85;
wire mux_o_86;
wire mux_o_87;
wire mux_o_88;
wire mux_o_90;
wire mux_o_91;
wire mux_o_92;
wire mux_o_93;
wire mux_o_94;
wire mux_o_95;
wire mux_o_97;
wire mux_o_98;
wire mux_o_99;
wire mux_o_101;
wire mux_o_102;
wire mux_o_104;
wire mux_o_105;
wire mux_o_106;
wire mux_o_107;
wire mux_o_108;
wire mux_o_109;
wire mux_o_110;
wire mux_o_111;
wire mux_o_112;
wire mux_o_113;
wire mux_o_114;
wire mux_o_115;
wire mux_o_116;
wire mux_o_117;
wire mux_o_118;
wire mux_o_119;
wire mux_o_120;
wire mux_o_121;
wire mux_o_122;
wire mux_o_123;
wire mux_o_124;
wire mux_o_125;
wire mux_o_126;
wire mux_o_127;
wire mux_o_128;
wire mux_o_129;
wire mux_o_130;
wire mux_o_131;
wire mux_o_132;
wire mux_o_133;
wire mux_o_134;
wire mux_o_135;
wire mux_o_136;
wire mux_o_137;
wire mux_o_138;
wire mux_o_139;
wire mux_o_140;
wire mux_o_142;
wire mux_o_143;
wire mux_o_144;
wire mux_o_145;
wire mux_o_146;
wire mux_o_147;
wire mux_o_149;
wire mux_o_150;
wire mux_o_151;
wire mux_o_153;
wire mux_o_154;
wire mux_o_156;
wire mux_o_157;
wire mux_o_158;
wire mux_o_159;
wire mux_o_160;
wire mux_o_161;
wire mux_o_162;
wire mux_o_163;
wire mux_o_164;
wire mux_o_165;
wire mux_o_166;
wire mux_o_167;
wire mux_o_168;
wire mux_o_169;
wire mux_o_170;
wire mux_o_171;
wire mux_o_172;
wire mux_o_173;
wire mux_o_174;
wire mux_o_175;
wire mux_o_176;
wire mux_o_177;
wire mux_o_178;
wire mux_o_179;
wire mux_o_180;
wire mux_o_181;
wire mux_o_182;
wire mux_o_183;
wire mux_o_184;
wire mux_o_185;
wire mux_o_186;
wire mux_o_187;
wire mux_o_188;
wire mux_o_189;
wire mux_o_190;
wire mux_o_191;
wire mux_o_192;
wire mux_o_194;
wire mux_o_195;
wire mux_o_196;
wire mux_o_197;
wire mux_o_198;
wire mux_o_199;
wire mux_o_201;
wire mux_o_202;
wire mux_o_203;
wire mux_o_205;
wire mux_o_206;
wire mux_o_208;
wire mux_o_209;
wire mux_o_210;
wire mux_o_211;
wire mux_o_212;
wire mux_o_213;
wire mux_o_214;
wire mux_o_215;
wire mux_o_216;
wire mux_o_217;
wire mux_o_218;
wire mux_o_219;
wire mux_o_220;
wire mux_o_221;
wire mux_o_222;
wire mux_o_223;
wire mux_o_224;
wire mux_o_225;
wire mux_o_226;
wire mux_o_227;
wire mux_o_228;
wire mux_o_229;
wire mux_o_230;
wire mux_o_231;
wire mux_o_232;
wire mux_o_233;
wire mux_o_234;
wire mux_o_235;
wire mux_o_236;
wire mux_o_237;
wire mux_o_238;
wire mux_o_239;
wire mux_o_240;
wire mux_o_241;
wire mux_o_242;
wire mux_o_243;
wire mux_o_244;
wire mux_o_246;
wire mux_o_247;
wire mux_o_248;
wire mux_o_249;
wire mux_o_250;
wire mux_o_251;
wire mux_o_253;
wire mux_o_254;
wire mux_o_255;
wire mux_o_257;
wire mux_o_258;
wire mux_o_260;
wire mux_o_261;
wire mux_o_262;
wire mux_o_263;
wire mux_o_264;
wire mux_o_265;
wire mux_o_266;
wire mux_o_267;
wire mux_o_268;
wire mux_o_269;
wire mux_o_270;
wire mux_o_271;
wire mux_o_272;
wire mux_o_273;
wire mux_o_274;
wire mux_o_275;
wire mux_o_276;
wire mux_o_277;
wire mux_o_278;
wire mux_o_279;
wire mux_o_280;
wire mux_o_281;
wire mux_o_282;
wire mux_o_283;
wire mux_o_284;
wire mux_o_285;
wire mux_o_286;
wire mux_o_287;
wire mux_o_288;
wire mux_o_289;
wire mux_o_290;
wire mux_o_291;
wire mux_o_292;
wire mux_o_293;
wire mux_o_294;
wire mux_o_295;
wire mux_o_296;
wire mux_o_298;
wire mux_o_299;
wire mux_o_300;
wire mux_o_301;
wire mux_o_302;
wire mux_o_303;
wire mux_o_305;
wire mux_o_306;
wire mux_o_307;
wire mux_o_309;
wire mux_o_310;
wire mux_o_312;
wire mux_o_313;
wire mux_o_314;
wire mux_o_315;
wire mux_o_316;
wire mux_o_317;
wire mux_o_318;
wire mux_o_319;
wire mux_o_320;
wire mux_o_321;
wire mux_o_322;
wire mux_o_323;
wire mux_o_324;
wire mux_o_325;
wire mux_o_326;
wire mux_o_327;
wire mux_o_328;
wire mux_o_329;
wire mux_o_330;
wire mux_o_331;
wire mux_o_332;
wire mux_o_333;
wire mux_o_334;
wire mux_o_335;
wire mux_o_336;
wire mux_o_337;
wire mux_o_338;
wire mux_o_339;
wire mux_o_340;
wire mux_o_341;
wire mux_o_342;
wire mux_o_343;
wire mux_o_344;
wire mux_o_345;
wire mux_o_346;
wire mux_o_347;
wire mux_o_348;
wire mux_o_350;
wire mux_o_351;
wire mux_o_352;
wire mux_o_353;
wire mux_o_354;
wire mux_o_355;
wire mux_o_357;
wire mux_o_358;
wire mux_o_359;
wire mux_o_361;
wire mux_o_362;
wire mux_o_364;
wire mux_o_365;
wire mux_o_366;
wire mux_o_367;
wire mux_o_368;
wire mux_o_369;
wire mux_o_370;
wire mux_o_371;
wire mux_o_372;
wire mux_o_373;
wire mux_o_374;
wire mux_o_375;
wire mux_o_376;
wire mux_o_377;
wire mux_o_378;
wire mux_o_379;
wire mux_o_380;
wire mux_o_381;
wire mux_o_382;
wire mux_o_383;
wire mux_o_384;
wire mux_o_385;
wire mux_o_386;
wire mux_o_387;
wire mux_o_388;
wire mux_o_389;
wire mux_o_390;
wire mux_o_391;
wire mux_o_392;
wire mux_o_393;
wire mux_o_394;
wire mux_o_395;
wire mux_o_396;
wire mux_o_397;
wire mux_o_398;
wire mux_o_399;
wire mux_o_400;
wire mux_o_402;
wire mux_o_403;
wire mux_o_404;
wire mux_o_405;
wire mux_o_406;
wire mux_o_407;
wire mux_o_409;
wire mux_o_410;
wire mux_o_411;
wire mux_o_413;
wire mux_o_414;

INV inv_inst_0 (.I(wad[4]), .O(wad4_inv));

INV inv_inst_1 (.I(wad[5]), .O(wad5_inv));

INV inv_inst_2 (.I(wad[6]), .O(wad6_inv));

INV inv_inst_3 (.I(wad[7]), .O(wad7_inv));

INV inv_inst_4 (.I(wad[8]), .O(wad8_inv));

INV inv_inst_5 (.I(wad[9]), .O(wad9_inv));

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_0.INIT = 16'h8000;
LUT4 lut_inst_1 (
  .F(lut_f_1),
  .I0(lut_f_0),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_1.INIT = 16'h8000;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_2.INIT = 16'h8000;
LUT4 lut_inst_3 (
  .F(lut_f_3),
  .I0(lut_f_2),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_3.INIT = 16'h8000;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_4.INIT = 16'h8000;
LUT4 lut_inst_5 (
  .F(lut_f_5),
  .I0(lut_f_4),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_5.INIT = 16'h8000;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_6.INIT = 16'h8000;
LUT4 lut_inst_7 (
  .F(lut_f_7),
  .I0(lut_f_6),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_7.INIT = 16'h8000;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_8.INIT = 16'h8000;
LUT4 lut_inst_9 (
  .F(lut_f_9),
  .I0(lut_f_8),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_9.INIT = 16'h8000;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_10.INIT = 16'h8000;
LUT4 lut_inst_11 (
  .F(lut_f_11),
  .I0(lut_f_10),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_11.INIT = 16'h8000;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_12.INIT = 16'h8000;
LUT4 lut_inst_13 (
  .F(lut_f_13),
  .I0(lut_f_12),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_13.INIT = 16'h8000;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_14.INIT = 16'h8000;
LUT4 lut_inst_15 (
  .F(lut_f_15),
  .I0(lut_f_14),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_15.INIT = 16'h8000;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_16.INIT = 16'h8000;
LUT4 lut_inst_17 (
  .F(lut_f_17),
  .I0(lut_f_16),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_17.INIT = 16'h8000;
LUT4 lut_inst_18 (
  .F(lut_f_18),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_18.INIT = 16'h8000;
LUT4 lut_inst_19 (
  .F(lut_f_19),
  .I0(lut_f_18),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_19.INIT = 16'h8000;
LUT4 lut_inst_20 (
  .F(lut_f_20),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_20.INIT = 16'h8000;
LUT4 lut_inst_21 (
  .F(lut_f_21),
  .I0(lut_f_20),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_21.INIT = 16'h8000;
LUT4 lut_inst_22 (
  .F(lut_f_22),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_22.INIT = 16'h8000;
LUT4 lut_inst_23 (
  .F(lut_f_23),
  .I0(lut_f_22),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_23.INIT = 16'h8000;
LUT4 lut_inst_24 (
  .F(lut_f_24),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_24.INIT = 16'h8000;
LUT4 lut_inst_25 (
  .F(lut_f_25),
  .I0(lut_f_24),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_25.INIT = 16'h8000;
LUT4 lut_inst_26 (
  .F(lut_f_26),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_26.INIT = 16'h8000;
LUT4 lut_inst_27 (
  .F(lut_f_27),
  .I0(lut_f_26),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_27.INIT = 16'h8000;
LUT4 lut_inst_28 (
  .F(lut_f_28),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_28.INIT = 16'h8000;
LUT4 lut_inst_29 (
  .F(lut_f_29),
  .I0(lut_f_28),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_29.INIT = 16'h8000;
LUT4 lut_inst_30 (
  .F(lut_f_30),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_30.INIT = 16'h8000;
LUT4 lut_inst_31 (
  .F(lut_f_31),
  .I0(lut_f_30),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad9_inv)
);
defparam lut_inst_31.INIT = 16'h8000;
LUT4 lut_inst_32 (
  .F(lut_f_32),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_32.INIT = 16'h8000;
LUT4 lut_inst_33 (
  .F(lut_f_33),
  .I0(lut_f_32),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_33.INIT = 16'h8000;
LUT4 lut_inst_34 (
  .F(lut_f_34),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_34.INIT = 16'h8000;
LUT4 lut_inst_35 (
  .F(lut_f_35),
  .I0(lut_f_34),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_35.INIT = 16'h8000;
LUT4 lut_inst_36 (
  .F(lut_f_36),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_36.INIT = 16'h8000;
LUT4 lut_inst_37 (
  .F(lut_f_37),
  .I0(lut_f_36),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_37.INIT = 16'h8000;
LUT4 lut_inst_38 (
  .F(lut_f_38),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_38.INIT = 16'h8000;
LUT4 lut_inst_39 (
  .F(lut_f_39),
  .I0(lut_f_38),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_39.INIT = 16'h8000;
LUT4 lut_inst_40 (
  .F(lut_f_40),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_40.INIT = 16'h8000;
LUT4 lut_inst_41 (
  .F(lut_f_41),
  .I0(lut_f_40),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_41.INIT = 16'h8000;
LUT4 lut_inst_42 (
  .F(lut_f_42),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_42.INIT = 16'h8000;
LUT4 lut_inst_43 (
  .F(lut_f_43),
  .I0(lut_f_42),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_43.INIT = 16'h8000;
LUT4 lut_inst_44 (
  .F(lut_f_44),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_44.INIT = 16'h8000;
LUT4 lut_inst_45 (
  .F(lut_f_45),
  .I0(lut_f_44),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_45.INIT = 16'h8000;
LUT4 lut_inst_46 (
  .F(lut_f_46),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_46.INIT = 16'h8000;
LUT4 lut_inst_47 (
  .F(lut_f_47),
  .I0(lut_f_46),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_47.INIT = 16'h8000;
LUT4 lut_inst_48 (
  .F(lut_f_48),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_48.INIT = 16'h8000;
LUT4 lut_inst_49 (
  .F(lut_f_49),
  .I0(lut_f_48),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_49.INIT = 16'h8000;
LUT4 lut_inst_50 (
  .F(lut_f_50),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_50.INIT = 16'h8000;
LUT4 lut_inst_51 (
  .F(lut_f_51),
  .I0(lut_f_50),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_51.INIT = 16'h8000;
LUT4 lut_inst_52 (
  .F(lut_f_52),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_52.INIT = 16'h8000;
LUT4 lut_inst_53 (
  .F(lut_f_53),
  .I0(lut_f_52),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_53.INIT = 16'h8000;
LUT4 lut_inst_54 (
  .F(lut_f_54),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_54.INIT = 16'h8000;
LUT4 lut_inst_55 (
  .F(lut_f_55),
  .I0(lut_f_54),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_55.INIT = 16'h8000;
LUT4 lut_inst_56 (
  .F(lut_f_56),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_56.INIT = 16'h8000;
LUT4 lut_inst_57 (
  .F(lut_f_57),
  .I0(lut_f_56),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_57.INIT = 16'h8000;
LUT4 lut_inst_58 (
  .F(lut_f_58),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_58.INIT = 16'h8000;
LUT4 lut_inst_59 (
  .F(lut_f_59),
  .I0(lut_f_58),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_59.INIT = 16'h8000;
LUT4 lut_inst_60 (
  .F(lut_f_60),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_60.INIT = 16'h8000;
LUT4 lut_inst_61 (
  .F(lut_f_61),
  .I0(lut_f_60),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_61.INIT = 16'h8000;
LUT4 lut_inst_62 (
  .F(lut_f_62),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_62.INIT = 16'h8000;
LUT4 lut_inst_63 (
  .F(lut_f_63),
  .I0(lut_f_62),
  .I1(wad[7]),
  .I2(wad[8]),
  .I3(wad9_inv)
);
defparam lut_inst_63.INIT = 16'h8000;
LUT4 lut_inst_64 (
  .F(lut_f_64),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_64.INIT = 16'h8000;
LUT4 lut_inst_65 (
  .F(lut_f_65),
  .I0(lut_f_64),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_65.INIT = 16'h8000;
LUT4 lut_inst_66 (
  .F(lut_f_66),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_66.INIT = 16'h8000;
LUT4 lut_inst_67 (
  .F(lut_f_67),
  .I0(lut_f_66),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_67.INIT = 16'h8000;
LUT4 lut_inst_68 (
  .F(lut_f_68),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_68.INIT = 16'h8000;
LUT4 lut_inst_69 (
  .F(lut_f_69),
  .I0(lut_f_68),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_69.INIT = 16'h8000;
LUT4 lut_inst_70 (
  .F(lut_f_70),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_70.INIT = 16'h8000;
LUT4 lut_inst_71 (
  .F(lut_f_71),
  .I0(lut_f_70),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_71.INIT = 16'h8000;
LUT4 lut_inst_72 (
  .F(lut_f_72),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_72.INIT = 16'h8000;
LUT4 lut_inst_73 (
  .F(lut_f_73),
  .I0(lut_f_72),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_73.INIT = 16'h8000;
LUT4 lut_inst_74 (
  .F(lut_f_74),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_74.INIT = 16'h8000;
LUT4 lut_inst_75 (
  .F(lut_f_75),
  .I0(lut_f_74),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_75.INIT = 16'h8000;
LUT4 lut_inst_76 (
  .F(lut_f_76),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_76.INIT = 16'h8000;
LUT4 lut_inst_77 (
  .F(lut_f_77),
  .I0(lut_f_76),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_77.INIT = 16'h8000;
LUT4 lut_inst_78 (
  .F(lut_f_78),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_78.INIT = 16'h8000;
LUT4 lut_inst_79 (
  .F(lut_f_79),
  .I0(lut_f_78),
  .I1(wad7_inv),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_79.INIT = 16'h8000;
LUT4 lut_inst_80 (
  .F(lut_f_80),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_80.INIT = 16'h8000;
LUT4 lut_inst_81 (
  .F(lut_f_81),
  .I0(lut_f_80),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_81.INIT = 16'h8000;
LUT4 lut_inst_82 (
  .F(lut_f_82),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_82.INIT = 16'h8000;
LUT4 lut_inst_83 (
  .F(lut_f_83),
  .I0(lut_f_82),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_83.INIT = 16'h8000;
LUT4 lut_inst_84 (
  .F(lut_f_84),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_84.INIT = 16'h8000;
LUT4 lut_inst_85 (
  .F(lut_f_85),
  .I0(lut_f_84),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_85.INIT = 16'h8000;
LUT4 lut_inst_86 (
  .F(lut_f_86),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad6_inv)
);
defparam lut_inst_86.INIT = 16'h8000;
LUT4 lut_inst_87 (
  .F(lut_f_87),
  .I0(lut_f_86),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_87.INIT = 16'h8000;
LUT4 lut_inst_88 (
  .F(lut_f_88),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_88.INIT = 16'h8000;
LUT4 lut_inst_89 (
  .F(lut_f_89),
  .I0(lut_f_88),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_89.INIT = 16'h8000;
LUT4 lut_inst_90 (
  .F(lut_f_90),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad[6])
);
defparam lut_inst_90.INIT = 16'h8000;
LUT4 lut_inst_91 (
  .F(lut_f_91),
  .I0(lut_f_90),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_91.INIT = 16'h8000;
LUT4 lut_inst_92 (
  .F(lut_f_92),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_92.INIT = 16'h8000;
LUT4 lut_inst_93 (
  .F(lut_f_93),
  .I0(lut_f_92),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_93.INIT = 16'h8000;
LUT4 lut_inst_94 (
  .F(lut_f_94),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad[5]),
  .I3(wad[6])
);
defparam lut_inst_94.INIT = 16'h8000;
LUT4 lut_inst_95 (
  .F(lut_f_95),
  .I0(lut_f_94),
  .I1(wad[7]),
  .I2(wad8_inv),
  .I3(wad[9])
);
defparam lut_inst_95.INIT = 16'h8000;
LUT4 lut_inst_96 (
  .F(lut_f_96),
  .I0(wre),
  .I1(wad4_inv),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_96.INIT = 16'h8000;
LUT4 lut_inst_97 (
  .F(lut_f_97),
  .I0(lut_f_96),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad[9])
);
defparam lut_inst_97.INIT = 16'h8000;
LUT4 lut_inst_98 (
  .F(lut_f_98),
  .I0(wre),
  .I1(wad[4]),
  .I2(wad5_inv),
  .I3(wad6_inv)
);
defparam lut_inst_98.INIT = 16'h8000;
LUT4 lut_inst_99 (
  .F(lut_f_99),
  .I0(lut_f_98),
  .I1(wad7_inv),
  .I2(wad[8]),
  .I3(wad[9])
);
defparam lut_inst_99.INIT = 16'h8000;
RAM16SDP4 ram16sdp_inst_0 (
    .DO(ram16sdp_inst_0_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16sdp_inst_0.INIT_0 = 16'h0000;
defparam ram16sdp_inst_0.INIT_1 = 16'h0000;
defparam ram16sdp_inst_0.INIT_2 = 16'h0000;
defparam ram16sdp_inst_0.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_1 (
    .DO(ram16sdp_inst_1_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_1),
    .CLK(clk)
);

defparam ram16sdp_inst_1.INIT_0 = 16'h0000;
defparam ram16sdp_inst_1.INIT_1 = 16'h0000;
defparam ram16sdp_inst_1.INIT_2 = 16'h0000;
defparam ram16sdp_inst_1.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_2 (
    .DO(ram16sdp_inst_2_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_3),
    .CLK(clk)
);

defparam ram16sdp_inst_2.INIT_0 = 16'h0000;
defparam ram16sdp_inst_2.INIT_1 = 16'h0000;
defparam ram16sdp_inst_2.INIT_2 = 16'h0000;
defparam ram16sdp_inst_2.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_3 (
    .DO(ram16sdp_inst_3_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_3),
    .CLK(clk)
);

defparam ram16sdp_inst_3.INIT_0 = 16'h0000;
defparam ram16sdp_inst_3.INIT_1 = 16'h0000;
defparam ram16sdp_inst_3.INIT_2 = 16'h0000;
defparam ram16sdp_inst_3.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_4 (
    .DO(ram16sdp_inst_4_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_4.INIT_0 = 16'h0000;
defparam ram16sdp_inst_4.INIT_1 = 16'h0000;
defparam ram16sdp_inst_4.INIT_2 = 16'h0000;
defparam ram16sdp_inst_4.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_5 (
    .DO(ram16sdp_inst_5_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_5),
    .CLK(clk)
);

defparam ram16sdp_inst_5.INIT_0 = 16'h0000;
defparam ram16sdp_inst_5.INIT_1 = 16'h0000;
defparam ram16sdp_inst_5.INIT_2 = 16'h0000;
defparam ram16sdp_inst_5.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_6 (
    .DO(ram16sdp_inst_6_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_7),
    .CLK(clk)
);

defparam ram16sdp_inst_6.INIT_0 = 16'h0000;
defparam ram16sdp_inst_6.INIT_1 = 16'h0000;
defparam ram16sdp_inst_6.INIT_2 = 16'h0000;
defparam ram16sdp_inst_6.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_7 (
    .DO(ram16sdp_inst_7_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_7),
    .CLK(clk)
);

defparam ram16sdp_inst_7.INIT_0 = 16'h0000;
defparam ram16sdp_inst_7.INIT_1 = 16'h0000;
defparam ram16sdp_inst_7.INIT_2 = 16'h0000;
defparam ram16sdp_inst_7.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_8 (
    .DO(ram16sdp_inst_8_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_9),
    .CLK(clk)
);

defparam ram16sdp_inst_8.INIT_0 = 16'h0000;
defparam ram16sdp_inst_8.INIT_1 = 16'h0000;
defparam ram16sdp_inst_8.INIT_2 = 16'h0000;
defparam ram16sdp_inst_8.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_9 (
    .DO(ram16sdp_inst_9_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_9),
    .CLK(clk)
);

defparam ram16sdp_inst_9.INIT_0 = 16'h0000;
defparam ram16sdp_inst_9.INIT_1 = 16'h0000;
defparam ram16sdp_inst_9.INIT_2 = 16'h0000;
defparam ram16sdp_inst_9.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_10 (
    .DO(ram16sdp_inst_10_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_10.INIT_0 = 16'h0000;
defparam ram16sdp_inst_10.INIT_1 = 16'h0000;
defparam ram16sdp_inst_10.INIT_2 = 16'h0000;
defparam ram16sdp_inst_10.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_11 (
    .DO(ram16sdp_inst_11_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_11),
    .CLK(clk)
);

defparam ram16sdp_inst_11.INIT_0 = 16'h0000;
defparam ram16sdp_inst_11.INIT_1 = 16'h0000;
defparam ram16sdp_inst_11.INIT_2 = 16'h0000;
defparam ram16sdp_inst_11.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_12 (
    .DO(ram16sdp_inst_12_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_13),
    .CLK(clk)
);

defparam ram16sdp_inst_12.INIT_0 = 16'h0000;
defparam ram16sdp_inst_12.INIT_1 = 16'h0000;
defparam ram16sdp_inst_12.INIT_2 = 16'h0000;
defparam ram16sdp_inst_12.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_13 (
    .DO(ram16sdp_inst_13_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_13),
    .CLK(clk)
);

defparam ram16sdp_inst_13.INIT_0 = 16'h0000;
defparam ram16sdp_inst_13.INIT_1 = 16'h0000;
defparam ram16sdp_inst_13.INIT_2 = 16'h0000;
defparam ram16sdp_inst_13.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_14 (
    .DO(ram16sdp_inst_14_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_15),
    .CLK(clk)
);

defparam ram16sdp_inst_14.INIT_0 = 16'h0000;
defparam ram16sdp_inst_14.INIT_1 = 16'h0000;
defparam ram16sdp_inst_14.INIT_2 = 16'h0000;
defparam ram16sdp_inst_14.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_15 (
    .DO(ram16sdp_inst_15_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_15),
    .CLK(clk)
);

defparam ram16sdp_inst_15.INIT_0 = 16'h0000;
defparam ram16sdp_inst_15.INIT_1 = 16'h0000;
defparam ram16sdp_inst_15.INIT_2 = 16'h0000;
defparam ram16sdp_inst_15.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_16 (
    .DO(ram16sdp_inst_16_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_16.INIT_0 = 16'h0000;
defparam ram16sdp_inst_16.INIT_1 = 16'h0000;
defparam ram16sdp_inst_16.INIT_2 = 16'h0000;
defparam ram16sdp_inst_16.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_17 (
    .DO(ram16sdp_inst_17_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_17),
    .CLK(clk)
);

defparam ram16sdp_inst_17.INIT_0 = 16'h0000;
defparam ram16sdp_inst_17.INIT_1 = 16'h0000;
defparam ram16sdp_inst_17.INIT_2 = 16'h0000;
defparam ram16sdp_inst_17.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_18 (
    .DO(ram16sdp_inst_18_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_19),
    .CLK(clk)
);

defparam ram16sdp_inst_18.INIT_0 = 16'h0000;
defparam ram16sdp_inst_18.INIT_1 = 16'h0000;
defparam ram16sdp_inst_18.INIT_2 = 16'h0000;
defparam ram16sdp_inst_18.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_19 (
    .DO(ram16sdp_inst_19_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_19),
    .CLK(clk)
);

defparam ram16sdp_inst_19.INIT_0 = 16'h0000;
defparam ram16sdp_inst_19.INIT_1 = 16'h0000;
defparam ram16sdp_inst_19.INIT_2 = 16'h0000;
defparam ram16sdp_inst_19.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_20 (
    .DO(ram16sdp_inst_20_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_21),
    .CLK(clk)
);

defparam ram16sdp_inst_20.INIT_0 = 16'h0000;
defparam ram16sdp_inst_20.INIT_1 = 16'h0000;
defparam ram16sdp_inst_20.INIT_2 = 16'h0000;
defparam ram16sdp_inst_20.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_21 (
    .DO(ram16sdp_inst_21_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_21),
    .CLK(clk)
);

defparam ram16sdp_inst_21.INIT_0 = 16'h0000;
defparam ram16sdp_inst_21.INIT_1 = 16'h0000;
defparam ram16sdp_inst_21.INIT_2 = 16'h0000;
defparam ram16sdp_inst_21.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_22 (
    .DO(ram16sdp_inst_22_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_22.INIT_0 = 16'h0000;
defparam ram16sdp_inst_22.INIT_1 = 16'h0000;
defparam ram16sdp_inst_22.INIT_2 = 16'h0000;
defparam ram16sdp_inst_22.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_23 (
    .DO(ram16sdp_inst_23_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_23),
    .CLK(clk)
);

defparam ram16sdp_inst_23.INIT_0 = 16'h0000;
defparam ram16sdp_inst_23.INIT_1 = 16'h0000;
defparam ram16sdp_inst_23.INIT_2 = 16'h0000;
defparam ram16sdp_inst_23.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_24 (
    .DO(ram16sdp_inst_24_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_25),
    .CLK(clk)
);

defparam ram16sdp_inst_24.INIT_0 = 16'h0000;
defparam ram16sdp_inst_24.INIT_1 = 16'h0000;
defparam ram16sdp_inst_24.INIT_2 = 16'h0000;
defparam ram16sdp_inst_24.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_25 (
    .DO(ram16sdp_inst_25_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_25),
    .CLK(clk)
);

defparam ram16sdp_inst_25.INIT_0 = 16'h0000;
defparam ram16sdp_inst_25.INIT_1 = 16'h0000;
defparam ram16sdp_inst_25.INIT_2 = 16'h0000;
defparam ram16sdp_inst_25.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_26 (
    .DO(ram16sdp_inst_26_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_27),
    .CLK(clk)
);

defparam ram16sdp_inst_26.INIT_0 = 16'h0000;
defparam ram16sdp_inst_26.INIT_1 = 16'h0000;
defparam ram16sdp_inst_26.INIT_2 = 16'h0000;
defparam ram16sdp_inst_26.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_27 (
    .DO(ram16sdp_inst_27_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_27),
    .CLK(clk)
);

defparam ram16sdp_inst_27.INIT_0 = 16'h0000;
defparam ram16sdp_inst_27.INIT_1 = 16'h0000;
defparam ram16sdp_inst_27.INIT_2 = 16'h0000;
defparam ram16sdp_inst_27.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_28 (
    .DO(ram16sdp_inst_28_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_28.INIT_0 = 16'h0000;
defparam ram16sdp_inst_28.INIT_1 = 16'h0000;
defparam ram16sdp_inst_28.INIT_2 = 16'h0000;
defparam ram16sdp_inst_28.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_29 (
    .DO(ram16sdp_inst_29_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_29),
    .CLK(clk)
);

defparam ram16sdp_inst_29.INIT_0 = 16'h0000;
defparam ram16sdp_inst_29.INIT_1 = 16'h0000;
defparam ram16sdp_inst_29.INIT_2 = 16'h0000;
defparam ram16sdp_inst_29.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_30 (
    .DO(ram16sdp_inst_30_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_31),
    .CLK(clk)
);

defparam ram16sdp_inst_30.INIT_0 = 16'h0000;
defparam ram16sdp_inst_30.INIT_1 = 16'h0000;
defparam ram16sdp_inst_30.INIT_2 = 16'h0000;
defparam ram16sdp_inst_30.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_31 (
    .DO(ram16sdp_inst_31_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_31),
    .CLK(clk)
);

defparam ram16sdp_inst_31.INIT_0 = 16'h0000;
defparam ram16sdp_inst_31.INIT_1 = 16'h0000;
defparam ram16sdp_inst_31.INIT_2 = 16'h0000;
defparam ram16sdp_inst_31.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_32 (
    .DO(ram16sdp_inst_32_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_33),
    .CLK(clk)
);

defparam ram16sdp_inst_32.INIT_0 = 16'h0000;
defparam ram16sdp_inst_32.INIT_1 = 16'h0000;
defparam ram16sdp_inst_32.INIT_2 = 16'h0000;
defparam ram16sdp_inst_32.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_33 (
    .DO(ram16sdp_inst_33_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_33),
    .CLK(clk)
);

defparam ram16sdp_inst_33.INIT_0 = 16'h0000;
defparam ram16sdp_inst_33.INIT_1 = 16'h0000;
defparam ram16sdp_inst_33.INIT_2 = 16'h0000;
defparam ram16sdp_inst_33.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_34 (
    .DO(ram16sdp_inst_34_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_34.INIT_0 = 16'h0000;
defparam ram16sdp_inst_34.INIT_1 = 16'h0000;
defparam ram16sdp_inst_34.INIT_2 = 16'h0000;
defparam ram16sdp_inst_34.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_35 (
    .DO(ram16sdp_inst_35_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_35),
    .CLK(clk)
);

defparam ram16sdp_inst_35.INIT_0 = 16'h0000;
defparam ram16sdp_inst_35.INIT_1 = 16'h0000;
defparam ram16sdp_inst_35.INIT_2 = 16'h0000;
defparam ram16sdp_inst_35.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_36 (
    .DO(ram16sdp_inst_36_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_37),
    .CLK(clk)
);

defparam ram16sdp_inst_36.INIT_0 = 16'h0000;
defparam ram16sdp_inst_36.INIT_1 = 16'h0000;
defparam ram16sdp_inst_36.INIT_2 = 16'h0000;
defparam ram16sdp_inst_36.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_37 (
    .DO(ram16sdp_inst_37_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_37),
    .CLK(clk)
);

defparam ram16sdp_inst_37.INIT_0 = 16'h0000;
defparam ram16sdp_inst_37.INIT_1 = 16'h0000;
defparam ram16sdp_inst_37.INIT_2 = 16'h0000;
defparam ram16sdp_inst_37.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_38 (
    .DO(ram16sdp_inst_38_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_39),
    .CLK(clk)
);

defparam ram16sdp_inst_38.INIT_0 = 16'h0000;
defparam ram16sdp_inst_38.INIT_1 = 16'h0000;
defparam ram16sdp_inst_38.INIT_2 = 16'h0000;
defparam ram16sdp_inst_38.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_39 (
    .DO(ram16sdp_inst_39_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_39),
    .CLK(clk)
);

defparam ram16sdp_inst_39.INIT_0 = 16'h0000;
defparam ram16sdp_inst_39.INIT_1 = 16'h0000;
defparam ram16sdp_inst_39.INIT_2 = 16'h0000;
defparam ram16sdp_inst_39.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_40 (
    .DO(ram16sdp_inst_40_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_40.INIT_0 = 16'h0000;
defparam ram16sdp_inst_40.INIT_1 = 16'h0000;
defparam ram16sdp_inst_40.INIT_2 = 16'h0000;
defparam ram16sdp_inst_40.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_41 (
    .DO(ram16sdp_inst_41_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_41),
    .CLK(clk)
);

defparam ram16sdp_inst_41.INIT_0 = 16'h0000;
defparam ram16sdp_inst_41.INIT_1 = 16'h0000;
defparam ram16sdp_inst_41.INIT_2 = 16'h0000;
defparam ram16sdp_inst_41.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_42 (
    .DO(ram16sdp_inst_42_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_43),
    .CLK(clk)
);

defparam ram16sdp_inst_42.INIT_0 = 16'h0000;
defparam ram16sdp_inst_42.INIT_1 = 16'h0000;
defparam ram16sdp_inst_42.INIT_2 = 16'h0000;
defparam ram16sdp_inst_42.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_43 (
    .DO(ram16sdp_inst_43_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_43),
    .CLK(clk)
);

defparam ram16sdp_inst_43.INIT_0 = 16'h0000;
defparam ram16sdp_inst_43.INIT_1 = 16'h0000;
defparam ram16sdp_inst_43.INIT_2 = 16'h0000;
defparam ram16sdp_inst_43.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_44 (
    .DO(ram16sdp_inst_44_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_45),
    .CLK(clk)
);

defparam ram16sdp_inst_44.INIT_0 = 16'h0000;
defparam ram16sdp_inst_44.INIT_1 = 16'h0000;
defparam ram16sdp_inst_44.INIT_2 = 16'h0000;
defparam ram16sdp_inst_44.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_45 (
    .DO(ram16sdp_inst_45_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_45),
    .CLK(clk)
);

defparam ram16sdp_inst_45.INIT_0 = 16'h0000;
defparam ram16sdp_inst_45.INIT_1 = 16'h0000;
defparam ram16sdp_inst_45.INIT_2 = 16'h0000;
defparam ram16sdp_inst_45.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_46 (
    .DO(ram16sdp_inst_46_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_46.INIT_0 = 16'h0000;
defparam ram16sdp_inst_46.INIT_1 = 16'h0000;
defparam ram16sdp_inst_46.INIT_2 = 16'h0000;
defparam ram16sdp_inst_46.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_47 (
    .DO(ram16sdp_inst_47_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_47),
    .CLK(clk)
);

defparam ram16sdp_inst_47.INIT_0 = 16'h0000;
defparam ram16sdp_inst_47.INIT_1 = 16'h0000;
defparam ram16sdp_inst_47.INIT_2 = 16'h0000;
defparam ram16sdp_inst_47.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_48 (
    .DO(ram16sdp_inst_48_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_49),
    .CLK(clk)
);

defparam ram16sdp_inst_48.INIT_0 = 16'h0000;
defparam ram16sdp_inst_48.INIT_1 = 16'h0000;
defparam ram16sdp_inst_48.INIT_2 = 16'h0000;
defparam ram16sdp_inst_48.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_49 (
    .DO(ram16sdp_inst_49_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_49),
    .CLK(clk)
);

defparam ram16sdp_inst_49.INIT_0 = 16'h0000;
defparam ram16sdp_inst_49.INIT_1 = 16'h0000;
defparam ram16sdp_inst_49.INIT_2 = 16'h0000;
defparam ram16sdp_inst_49.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_50 (
    .DO(ram16sdp_inst_50_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_51),
    .CLK(clk)
);

defparam ram16sdp_inst_50.INIT_0 = 16'h0000;
defparam ram16sdp_inst_50.INIT_1 = 16'h0000;
defparam ram16sdp_inst_50.INIT_2 = 16'h0000;
defparam ram16sdp_inst_50.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_51 (
    .DO(ram16sdp_inst_51_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_51),
    .CLK(clk)
);

defparam ram16sdp_inst_51.INIT_0 = 16'h0000;
defparam ram16sdp_inst_51.INIT_1 = 16'h0000;
defparam ram16sdp_inst_51.INIT_2 = 16'h0000;
defparam ram16sdp_inst_51.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_52 (
    .DO(ram16sdp_inst_52_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_52.INIT_0 = 16'h0000;
defparam ram16sdp_inst_52.INIT_1 = 16'h0000;
defparam ram16sdp_inst_52.INIT_2 = 16'h0000;
defparam ram16sdp_inst_52.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_53 (
    .DO(ram16sdp_inst_53_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_53),
    .CLK(clk)
);

defparam ram16sdp_inst_53.INIT_0 = 16'h0000;
defparam ram16sdp_inst_53.INIT_1 = 16'h0000;
defparam ram16sdp_inst_53.INIT_2 = 16'h0000;
defparam ram16sdp_inst_53.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_54 (
    .DO(ram16sdp_inst_54_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_55),
    .CLK(clk)
);

defparam ram16sdp_inst_54.INIT_0 = 16'h0000;
defparam ram16sdp_inst_54.INIT_1 = 16'h0000;
defparam ram16sdp_inst_54.INIT_2 = 16'h0000;
defparam ram16sdp_inst_54.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_55 (
    .DO(ram16sdp_inst_55_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_55),
    .CLK(clk)
);

defparam ram16sdp_inst_55.INIT_0 = 16'h0000;
defparam ram16sdp_inst_55.INIT_1 = 16'h0000;
defparam ram16sdp_inst_55.INIT_2 = 16'h0000;
defparam ram16sdp_inst_55.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_56 (
    .DO(ram16sdp_inst_56_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_57),
    .CLK(clk)
);

defparam ram16sdp_inst_56.INIT_0 = 16'h0000;
defparam ram16sdp_inst_56.INIT_1 = 16'h0000;
defparam ram16sdp_inst_56.INIT_2 = 16'h0000;
defparam ram16sdp_inst_56.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_57 (
    .DO(ram16sdp_inst_57_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_57),
    .CLK(clk)
);

defparam ram16sdp_inst_57.INIT_0 = 16'h0000;
defparam ram16sdp_inst_57.INIT_1 = 16'h0000;
defparam ram16sdp_inst_57.INIT_2 = 16'h0000;
defparam ram16sdp_inst_57.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_58 (
    .DO(ram16sdp_inst_58_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_58.INIT_0 = 16'h0000;
defparam ram16sdp_inst_58.INIT_1 = 16'h0000;
defparam ram16sdp_inst_58.INIT_2 = 16'h0000;
defparam ram16sdp_inst_58.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_59 (
    .DO(ram16sdp_inst_59_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_59),
    .CLK(clk)
);

defparam ram16sdp_inst_59.INIT_0 = 16'h0000;
defparam ram16sdp_inst_59.INIT_1 = 16'h0000;
defparam ram16sdp_inst_59.INIT_2 = 16'h0000;
defparam ram16sdp_inst_59.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_60 (
    .DO(ram16sdp_inst_60_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_61),
    .CLK(clk)
);

defparam ram16sdp_inst_60.INIT_0 = 16'h0000;
defparam ram16sdp_inst_60.INIT_1 = 16'h0000;
defparam ram16sdp_inst_60.INIT_2 = 16'h0000;
defparam ram16sdp_inst_60.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_61 (
    .DO(ram16sdp_inst_61_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_61),
    .CLK(clk)
);

defparam ram16sdp_inst_61.INIT_0 = 16'h0000;
defparam ram16sdp_inst_61.INIT_1 = 16'h0000;
defparam ram16sdp_inst_61.INIT_2 = 16'h0000;
defparam ram16sdp_inst_61.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_62 (
    .DO(ram16sdp_inst_62_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_63),
    .CLK(clk)
);

defparam ram16sdp_inst_62.INIT_0 = 16'h0000;
defparam ram16sdp_inst_62.INIT_1 = 16'h0000;
defparam ram16sdp_inst_62.INIT_2 = 16'h0000;
defparam ram16sdp_inst_62.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_63 (
    .DO(ram16sdp_inst_63_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_63),
    .CLK(clk)
);

defparam ram16sdp_inst_63.INIT_0 = 16'h0000;
defparam ram16sdp_inst_63.INIT_1 = 16'h0000;
defparam ram16sdp_inst_63.INIT_2 = 16'h0000;
defparam ram16sdp_inst_63.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_64 (
    .DO(ram16sdp_inst_64_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_64.INIT_0 = 16'h0000;
defparam ram16sdp_inst_64.INIT_1 = 16'h0000;
defparam ram16sdp_inst_64.INIT_2 = 16'h0000;
defparam ram16sdp_inst_64.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_65 (
    .DO(ram16sdp_inst_65_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_65),
    .CLK(clk)
);

defparam ram16sdp_inst_65.INIT_0 = 16'h0000;
defparam ram16sdp_inst_65.INIT_1 = 16'h0000;
defparam ram16sdp_inst_65.INIT_2 = 16'h0000;
defparam ram16sdp_inst_65.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_66 (
    .DO(ram16sdp_inst_66_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_67),
    .CLK(clk)
);

defparam ram16sdp_inst_66.INIT_0 = 16'h0000;
defparam ram16sdp_inst_66.INIT_1 = 16'h0000;
defparam ram16sdp_inst_66.INIT_2 = 16'h0000;
defparam ram16sdp_inst_66.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_67 (
    .DO(ram16sdp_inst_67_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_67),
    .CLK(clk)
);

defparam ram16sdp_inst_67.INIT_0 = 16'h0000;
defparam ram16sdp_inst_67.INIT_1 = 16'h0000;
defparam ram16sdp_inst_67.INIT_2 = 16'h0000;
defparam ram16sdp_inst_67.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_68 (
    .DO(ram16sdp_inst_68_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_69),
    .CLK(clk)
);

defparam ram16sdp_inst_68.INIT_0 = 16'h0000;
defparam ram16sdp_inst_68.INIT_1 = 16'h0000;
defparam ram16sdp_inst_68.INIT_2 = 16'h0000;
defparam ram16sdp_inst_68.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_69 (
    .DO(ram16sdp_inst_69_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_69),
    .CLK(clk)
);

defparam ram16sdp_inst_69.INIT_0 = 16'h0000;
defparam ram16sdp_inst_69.INIT_1 = 16'h0000;
defparam ram16sdp_inst_69.INIT_2 = 16'h0000;
defparam ram16sdp_inst_69.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_70 (
    .DO(ram16sdp_inst_70_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_70.INIT_0 = 16'h0000;
defparam ram16sdp_inst_70.INIT_1 = 16'h0000;
defparam ram16sdp_inst_70.INIT_2 = 16'h0000;
defparam ram16sdp_inst_70.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_71 (
    .DO(ram16sdp_inst_71_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_71),
    .CLK(clk)
);

defparam ram16sdp_inst_71.INIT_0 = 16'h0000;
defparam ram16sdp_inst_71.INIT_1 = 16'h0000;
defparam ram16sdp_inst_71.INIT_2 = 16'h0000;
defparam ram16sdp_inst_71.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_72 (
    .DO(ram16sdp_inst_72_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_73),
    .CLK(clk)
);

defparam ram16sdp_inst_72.INIT_0 = 16'h0000;
defparam ram16sdp_inst_72.INIT_1 = 16'h0000;
defparam ram16sdp_inst_72.INIT_2 = 16'h0000;
defparam ram16sdp_inst_72.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_73 (
    .DO(ram16sdp_inst_73_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_73),
    .CLK(clk)
);

defparam ram16sdp_inst_73.INIT_0 = 16'h0000;
defparam ram16sdp_inst_73.INIT_1 = 16'h0000;
defparam ram16sdp_inst_73.INIT_2 = 16'h0000;
defparam ram16sdp_inst_73.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_74 (
    .DO(ram16sdp_inst_74_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_75),
    .CLK(clk)
);

defparam ram16sdp_inst_74.INIT_0 = 16'h0000;
defparam ram16sdp_inst_74.INIT_1 = 16'h0000;
defparam ram16sdp_inst_74.INIT_2 = 16'h0000;
defparam ram16sdp_inst_74.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_75 (
    .DO(ram16sdp_inst_75_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_75),
    .CLK(clk)
);

defparam ram16sdp_inst_75.INIT_0 = 16'h0000;
defparam ram16sdp_inst_75.INIT_1 = 16'h0000;
defparam ram16sdp_inst_75.INIT_2 = 16'h0000;
defparam ram16sdp_inst_75.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_76 (
    .DO(ram16sdp_inst_76_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_76.INIT_0 = 16'h0000;
defparam ram16sdp_inst_76.INIT_1 = 16'h0000;
defparam ram16sdp_inst_76.INIT_2 = 16'h0000;
defparam ram16sdp_inst_76.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_77 (
    .DO(ram16sdp_inst_77_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_77),
    .CLK(clk)
);

defparam ram16sdp_inst_77.INIT_0 = 16'h0000;
defparam ram16sdp_inst_77.INIT_1 = 16'h0000;
defparam ram16sdp_inst_77.INIT_2 = 16'h0000;
defparam ram16sdp_inst_77.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_78 (
    .DO(ram16sdp_inst_78_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_79),
    .CLK(clk)
);

defparam ram16sdp_inst_78.INIT_0 = 16'h0000;
defparam ram16sdp_inst_78.INIT_1 = 16'h0000;
defparam ram16sdp_inst_78.INIT_2 = 16'h0000;
defparam ram16sdp_inst_78.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_79 (
    .DO(ram16sdp_inst_79_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_79),
    .CLK(clk)
);

defparam ram16sdp_inst_79.INIT_0 = 16'h0000;
defparam ram16sdp_inst_79.INIT_1 = 16'h0000;
defparam ram16sdp_inst_79.INIT_2 = 16'h0000;
defparam ram16sdp_inst_79.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_80 (
    .DO(ram16sdp_inst_80_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_81),
    .CLK(clk)
);

defparam ram16sdp_inst_80.INIT_0 = 16'h0000;
defparam ram16sdp_inst_80.INIT_1 = 16'h0000;
defparam ram16sdp_inst_80.INIT_2 = 16'h0000;
defparam ram16sdp_inst_80.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_81 (
    .DO(ram16sdp_inst_81_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_81),
    .CLK(clk)
);

defparam ram16sdp_inst_81.INIT_0 = 16'h0000;
defparam ram16sdp_inst_81.INIT_1 = 16'h0000;
defparam ram16sdp_inst_81.INIT_2 = 16'h0000;
defparam ram16sdp_inst_81.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_82 (
    .DO(ram16sdp_inst_82_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_82.INIT_0 = 16'h0000;
defparam ram16sdp_inst_82.INIT_1 = 16'h0000;
defparam ram16sdp_inst_82.INIT_2 = 16'h0000;
defparam ram16sdp_inst_82.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_83 (
    .DO(ram16sdp_inst_83_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_83),
    .CLK(clk)
);

defparam ram16sdp_inst_83.INIT_0 = 16'h0000;
defparam ram16sdp_inst_83.INIT_1 = 16'h0000;
defparam ram16sdp_inst_83.INIT_2 = 16'h0000;
defparam ram16sdp_inst_83.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_84 (
    .DO(ram16sdp_inst_84_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_85),
    .CLK(clk)
);

defparam ram16sdp_inst_84.INIT_0 = 16'h0000;
defparam ram16sdp_inst_84.INIT_1 = 16'h0000;
defparam ram16sdp_inst_84.INIT_2 = 16'h0000;
defparam ram16sdp_inst_84.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_85 (
    .DO(ram16sdp_inst_85_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_85),
    .CLK(clk)
);

defparam ram16sdp_inst_85.INIT_0 = 16'h0000;
defparam ram16sdp_inst_85.INIT_1 = 16'h0000;
defparam ram16sdp_inst_85.INIT_2 = 16'h0000;
defparam ram16sdp_inst_85.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_86 (
    .DO(ram16sdp_inst_86_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_87),
    .CLK(clk)
);

defparam ram16sdp_inst_86.INIT_0 = 16'h0000;
defparam ram16sdp_inst_86.INIT_1 = 16'h0000;
defparam ram16sdp_inst_86.INIT_2 = 16'h0000;
defparam ram16sdp_inst_86.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_87 (
    .DO(ram16sdp_inst_87_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_87),
    .CLK(clk)
);

defparam ram16sdp_inst_87.INIT_0 = 16'h0000;
defparam ram16sdp_inst_87.INIT_1 = 16'h0000;
defparam ram16sdp_inst_87.INIT_2 = 16'h0000;
defparam ram16sdp_inst_87.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_88 (
    .DO(ram16sdp_inst_88_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_88.INIT_0 = 16'h0000;
defparam ram16sdp_inst_88.INIT_1 = 16'h0000;
defparam ram16sdp_inst_88.INIT_2 = 16'h0000;
defparam ram16sdp_inst_88.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_89 (
    .DO(ram16sdp_inst_89_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_89),
    .CLK(clk)
);

defparam ram16sdp_inst_89.INIT_0 = 16'h0000;
defparam ram16sdp_inst_89.INIT_1 = 16'h0000;
defparam ram16sdp_inst_89.INIT_2 = 16'h0000;
defparam ram16sdp_inst_89.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_90 (
    .DO(ram16sdp_inst_90_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_91),
    .CLK(clk)
);

defparam ram16sdp_inst_90.INIT_0 = 16'h0000;
defparam ram16sdp_inst_90.INIT_1 = 16'h0000;
defparam ram16sdp_inst_90.INIT_2 = 16'h0000;
defparam ram16sdp_inst_90.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_91 (
    .DO(ram16sdp_inst_91_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_91),
    .CLK(clk)
);

defparam ram16sdp_inst_91.INIT_0 = 16'h0000;
defparam ram16sdp_inst_91.INIT_1 = 16'h0000;
defparam ram16sdp_inst_91.INIT_2 = 16'h0000;
defparam ram16sdp_inst_91.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_92 (
    .DO(ram16sdp_inst_92_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_93),
    .CLK(clk)
);

defparam ram16sdp_inst_92.INIT_0 = 16'h0000;
defparam ram16sdp_inst_92.INIT_1 = 16'h0000;
defparam ram16sdp_inst_92.INIT_2 = 16'h0000;
defparam ram16sdp_inst_92.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_93 (
    .DO(ram16sdp_inst_93_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_93),
    .CLK(clk)
);

defparam ram16sdp_inst_93.INIT_0 = 16'h0000;
defparam ram16sdp_inst_93.INIT_1 = 16'h0000;
defparam ram16sdp_inst_93.INIT_2 = 16'h0000;
defparam ram16sdp_inst_93.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_94 (
    .DO(ram16sdp_inst_94_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_94.INIT_0 = 16'h0000;
defparam ram16sdp_inst_94.INIT_1 = 16'h0000;
defparam ram16sdp_inst_94.INIT_2 = 16'h0000;
defparam ram16sdp_inst_94.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_95 (
    .DO(ram16sdp_inst_95_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_95),
    .CLK(clk)
);

defparam ram16sdp_inst_95.INIT_0 = 16'h0000;
defparam ram16sdp_inst_95.INIT_1 = 16'h0000;
defparam ram16sdp_inst_95.INIT_2 = 16'h0000;
defparam ram16sdp_inst_95.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_96 (
    .DO(ram16sdp_inst_96_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_97),
    .CLK(clk)
);

defparam ram16sdp_inst_96.INIT_0 = 16'h0000;
defparam ram16sdp_inst_96.INIT_1 = 16'h0000;
defparam ram16sdp_inst_96.INIT_2 = 16'h0000;
defparam ram16sdp_inst_96.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_97 (
    .DO(ram16sdp_inst_97_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_97),
    .CLK(clk)
);

defparam ram16sdp_inst_97.INIT_0 = 16'h0000;
defparam ram16sdp_inst_97.INIT_1 = 16'h0000;
defparam ram16sdp_inst_97.INIT_2 = 16'h0000;
defparam ram16sdp_inst_97.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_98 (
    .DO(ram16sdp_inst_98_dout[3:0]),
    .DI(di[3:0]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_99),
    .CLK(clk)
);

defparam ram16sdp_inst_98.INIT_0 = 16'h0000;
defparam ram16sdp_inst_98.INIT_1 = 16'h0000;
defparam ram16sdp_inst_98.INIT_2 = 16'h0000;
defparam ram16sdp_inst_98.INIT_3 = 16'h0000;

RAM16SDP4 ram16sdp_inst_99 (
    .DO(ram16sdp_inst_99_dout[7:4]),
    .DI(di[7:4]),
    .WAD(wad[3:0]),
    .RAD(rad[3:0]),
    .WRE(lut_f_99),
    .CLK(clk)
);

defparam ram16sdp_inst_99.INIT_0 = 16'h0000;
defparam ram16sdp_inst_99.INIT_1 = 16'h0000;
defparam ram16sdp_inst_99.INIT_2 = 16'h0000;
defparam ram16sdp_inst_99.INIT_3 = 16'h0000;

MUX2 mux_inst_0 (
  .O(mux_o_0),
  .I0(ram16sdp_inst_0_dout[0]),
  .I1(ram16sdp_inst_2_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_1 (
  .O(mux_o_1),
  .I0(ram16sdp_inst_4_dout[0]),
  .I1(ram16sdp_inst_6_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_2 (
  .O(mux_o_2),
  .I0(ram16sdp_inst_8_dout[0]),
  .I1(ram16sdp_inst_10_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_3 (
  .O(mux_o_3),
  .I0(ram16sdp_inst_12_dout[0]),
  .I1(ram16sdp_inst_14_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_4 (
  .O(mux_o_4),
  .I0(ram16sdp_inst_16_dout[0]),
  .I1(ram16sdp_inst_18_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_5 (
  .O(mux_o_5),
  .I0(ram16sdp_inst_20_dout[0]),
  .I1(ram16sdp_inst_22_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_6 (
  .O(mux_o_6),
  .I0(ram16sdp_inst_24_dout[0]),
  .I1(ram16sdp_inst_26_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_7 (
  .O(mux_o_7),
  .I0(ram16sdp_inst_28_dout[0]),
  .I1(ram16sdp_inst_30_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_8 (
  .O(mux_o_8),
  .I0(ram16sdp_inst_32_dout[0]),
  .I1(ram16sdp_inst_34_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_9 (
  .O(mux_o_9),
  .I0(ram16sdp_inst_36_dout[0]),
  .I1(ram16sdp_inst_38_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(ram16sdp_inst_40_dout[0]),
  .I1(ram16sdp_inst_42_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(ram16sdp_inst_44_dout[0]),
  .I1(ram16sdp_inst_46_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(ram16sdp_inst_48_dout[0]),
  .I1(ram16sdp_inst_50_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(ram16sdp_inst_52_dout[0]),
  .I1(ram16sdp_inst_54_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(ram16sdp_inst_56_dout[0]),
  .I1(ram16sdp_inst_58_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(ram16sdp_inst_60_dout[0]),
  .I1(ram16sdp_inst_62_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(ram16sdp_inst_64_dout[0]),
  .I1(ram16sdp_inst_66_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_17 (
  .O(mux_o_17),
  .I0(ram16sdp_inst_68_dout[0]),
  .I1(ram16sdp_inst_70_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(ram16sdp_inst_72_dout[0]),
  .I1(ram16sdp_inst_74_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_19 (
  .O(mux_o_19),
  .I0(ram16sdp_inst_76_dout[0]),
  .I1(ram16sdp_inst_78_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_20 (
  .O(mux_o_20),
  .I0(ram16sdp_inst_80_dout[0]),
  .I1(ram16sdp_inst_82_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_21 (
  .O(mux_o_21),
  .I0(ram16sdp_inst_84_dout[0]),
  .I1(ram16sdp_inst_86_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_22 (
  .O(mux_o_22),
  .I0(ram16sdp_inst_88_dout[0]),
  .I1(ram16sdp_inst_90_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_23 (
  .O(mux_o_23),
  .I0(ram16sdp_inst_92_dout[0]),
  .I1(ram16sdp_inst_94_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_24 (
  .O(mux_o_24),
  .I0(ram16sdp_inst_96_dout[0]),
  .I1(ram16sdp_inst_98_dout[0]),
  .S0(rad[4])
);
MUX2 mux_inst_25 (
  .O(mux_o_25),
  .I0(mux_o_0),
  .I1(mux_o_1),
  .S0(rad[5])
);
MUX2 mux_inst_26 (
  .O(mux_o_26),
  .I0(mux_o_2),
  .I1(mux_o_3),
  .S0(rad[5])
);
MUX2 mux_inst_27 (
  .O(mux_o_27),
  .I0(mux_o_4),
  .I1(mux_o_5),
  .S0(rad[5])
);
MUX2 mux_inst_28 (
  .O(mux_o_28),
  .I0(mux_o_6),
  .I1(mux_o_7),
  .S0(rad[5])
);
MUX2 mux_inst_29 (
  .O(mux_o_29),
  .I0(mux_o_8),
  .I1(mux_o_9),
  .S0(rad[5])
);
MUX2 mux_inst_30 (
  .O(mux_o_30),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(rad[5])
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(rad[5])
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(mux_o_14),
  .I1(mux_o_15),
  .S0(rad[5])
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(mux_o_16),
  .I1(mux_o_17),
  .S0(rad[5])
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(mux_o_18),
  .I1(mux_o_19),
  .S0(rad[5])
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(mux_o_20),
  .I1(mux_o_21),
  .S0(rad[5])
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(mux_o_22),
  .I1(mux_o_23),
  .S0(rad[5])
);
MUX2 mux_inst_38 (
  .O(mux_o_38),
  .I0(mux_o_25),
  .I1(mux_o_26),
  .S0(rad[6])
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_27),
  .I1(mux_o_28),
  .S0(rad[6])
);
MUX2 mux_inst_40 (
  .O(mux_o_40),
  .I0(mux_o_29),
  .I1(mux_o_30),
  .S0(rad[6])
);
MUX2 mux_inst_41 (
  .O(mux_o_41),
  .I0(mux_o_31),
  .I1(mux_o_32),
  .S0(rad[6])
);
MUX2 mux_inst_42 (
  .O(mux_o_42),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(rad[6])
);
MUX2 mux_inst_43 (
  .O(mux_o_43),
  .I0(mux_o_35),
  .I1(mux_o_36),
  .S0(rad[6])
);
MUX2 mux_inst_45 (
  .O(mux_o_45),
  .I0(mux_o_38),
  .I1(mux_o_39),
  .S0(rad[7])
);
MUX2 mux_inst_46 (
  .O(mux_o_46),
  .I0(mux_o_40),
  .I1(mux_o_41),
  .S0(rad[7])
);
MUX2 mux_inst_47 (
  .O(mux_o_47),
  .I0(mux_o_42),
  .I1(mux_o_43),
  .S0(rad[7])
);
MUX2 mux_inst_49 (
  .O(mux_o_49),
  .I0(mux_o_45),
  .I1(mux_o_46),
  .S0(rad[8])
);
MUX2 mux_inst_50 (
  .O(mux_o_50),
  .I0(mux_o_47),
  .I1(mux_o_24),
  .S0(rad[8])
);
MUX2 mux_inst_51 (
  .O(dout[0]),
  .I0(mux_o_49),
  .I1(mux_o_50),
  .S0(rad[9])
);
MUX2 mux_inst_52 (
  .O(mux_o_52),
  .I0(ram16sdp_inst_0_dout[1]),
  .I1(ram16sdp_inst_2_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_53 (
  .O(mux_o_53),
  .I0(ram16sdp_inst_4_dout[1]),
  .I1(ram16sdp_inst_6_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_54 (
  .O(mux_o_54),
  .I0(ram16sdp_inst_8_dout[1]),
  .I1(ram16sdp_inst_10_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_55 (
  .O(mux_o_55),
  .I0(ram16sdp_inst_12_dout[1]),
  .I1(ram16sdp_inst_14_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_56 (
  .O(mux_o_56),
  .I0(ram16sdp_inst_16_dout[1]),
  .I1(ram16sdp_inst_18_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_57 (
  .O(mux_o_57),
  .I0(ram16sdp_inst_20_dout[1]),
  .I1(ram16sdp_inst_22_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_58 (
  .O(mux_o_58),
  .I0(ram16sdp_inst_24_dout[1]),
  .I1(ram16sdp_inst_26_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_59 (
  .O(mux_o_59),
  .I0(ram16sdp_inst_28_dout[1]),
  .I1(ram16sdp_inst_30_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_60 (
  .O(mux_o_60),
  .I0(ram16sdp_inst_32_dout[1]),
  .I1(ram16sdp_inst_34_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_61 (
  .O(mux_o_61),
  .I0(ram16sdp_inst_36_dout[1]),
  .I1(ram16sdp_inst_38_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_62 (
  .O(mux_o_62),
  .I0(ram16sdp_inst_40_dout[1]),
  .I1(ram16sdp_inst_42_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_63 (
  .O(mux_o_63),
  .I0(ram16sdp_inst_44_dout[1]),
  .I1(ram16sdp_inst_46_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_64 (
  .O(mux_o_64),
  .I0(ram16sdp_inst_48_dout[1]),
  .I1(ram16sdp_inst_50_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_65 (
  .O(mux_o_65),
  .I0(ram16sdp_inst_52_dout[1]),
  .I1(ram16sdp_inst_54_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_66 (
  .O(mux_o_66),
  .I0(ram16sdp_inst_56_dout[1]),
  .I1(ram16sdp_inst_58_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_67 (
  .O(mux_o_67),
  .I0(ram16sdp_inst_60_dout[1]),
  .I1(ram16sdp_inst_62_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_68 (
  .O(mux_o_68),
  .I0(ram16sdp_inst_64_dout[1]),
  .I1(ram16sdp_inst_66_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_69 (
  .O(mux_o_69),
  .I0(ram16sdp_inst_68_dout[1]),
  .I1(ram16sdp_inst_70_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_70 (
  .O(mux_o_70),
  .I0(ram16sdp_inst_72_dout[1]),
  .I1(ram16sdp_inst_74_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_71 (
  .O(mux_o_71),
  .I0(ram16sdp_inst_76_dout[1]),
  .I1(ram16sdp_inst_78_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_72 (
  .O(mux_o_72),
  .I0(ram16sdp_inst_80_dout[1]),
  .I1(ram16sdp_inst_82_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_73 (
  .O(mux_o_73),
  .I0(ram16sdp_inst_84_dout[1]),
  .I1(ram16sdp_inst_86_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_74 (
  .O(mux_o_74),
  .I0(ram16sdp_inst_88_dout[1]),
  .I1(ram16sdp_inst_90_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_75 (
  .O(mux_o_75),
  .I0(ram16sdp_inst_92_dout[1]),
  .I1(ram16sdp_inst_94_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_76 (
  .O(mux_o_76),
  .I0(ram16sdp_inst_96_dout[1]),
  .I1(ram16sdp_inst_98_dout[1]),
  .S0(rad[4])
);
MUX2 mux_inst_77 (
  .O(mux_o_77),
  .I0(mux_o_52),
  .I1(mux_o_53),
  .S0(rad[5])
);
MUX2 mux_inst_78 (
  .O(mux_o_78),
  .I0(mux_o_54),
  .I1(mux_o_55),
  .S0(rad[5])
);
MUX2 mux_inst_79 (
  .O(mux_o_79),
  .I0(mux_o_56),
  .I1(mux_o_57),
  .S0(rad[5])
);
MUX2 mux_inst_80 (
  .O(mux_o_80),
  .I0(mux_o_58),
  .I1(mux_o_59),
  .S0(rad[5])
);
MUX2 mux_inst_81 (
  .O(mux_o_81),
  .I0(mux_o_60),
  .I1(mux_o_61),
  .S0(rad[5])
);
MUX2 mux_inst_82 (
  .O(mux_o_82),
  .I0(mux_o_62),
  .I1(mux_o_63),
  .S0(rad[5])
);
MUX2 mux_inst_83 (
  .O(mux_o_83),
  .I0(mux_o_64),
  .I1(mux_o_65),
  .S0(rad[5])
);
MUX2 mux_inst_84 (
  .O(mux_o_84),
  .I0(mux_o_66),
  .I1(mux_o_67),
  .S0(rad[5])
);
MUX2 mux_inst_85 (
  .O(mux_o_85),
  .I0(mux_o_68),
  .I1(mux_o_69),
  .S0(rad[5])
);
MUX2 mux_inst_86 (
  .O(mux_o_86),
  .I0(mux_o_70),
  .I1(mux_o_71),
  .S0(rad[5])
);
MUX2 mux_inst_87 (
  .O(mux_o_87),
  .I0(mux_o_72),
  .I1(mux_o_73),
  .S0(rad[5])
);
MUX2 mux_inst_88 (
  .O(mux_o_88),
  .I0(mux_o_74),
  .I1(mux_o_75),
  .S0(rad[5])
);
MUX2 mux_inst_90 (
  .O(mux_o_90),
  .I0(mux_o_77),
  .I1(mux_o_78),
  .S0(rad[6])
);
MUX2 mux_inst_91 (
  .O(mux_o_91),
  .I0(mux_o_79),
  .I1(mux_o_80),
  .S0(rad[6])
);
MUX2 mux_inst_92 (
  .O(mux_o_92),
  .I0(mux_o_81),
  .I1(mux_o_82),
  .S0(rad[6])
);
MUX2 mux_inst_93 (
  .O(mux_o_93),
  .I0(mux_o_83),
  .I1(mux_o_84),
  .S0(rad[6])
);
MUX2 mux_inst_94 (
  .O(mux_o_94),
  .I0(mux_o_85),
  .I1(mux_o_86),
  .S0(rad[6])
);
MUX2 mux_inst_95 (
  .O(mux_o_95),
  .I0(mux_o_87),
  .I1(mux_o_88),
  .S0(rad[6])
);
MUX2 mux_inst_97 (
  .O(mux_o_97),
  .I0(mux_o_90),
  .I1(mux_o_91),
  .S0(rad[7])
);
MUX2 mux_inst_98 (
  .O(mux_o_98),
  .I0(mux_o_92),
  .I1(mux_o_93),
  .S0(rad[7])
);
MUX2 mux_inst_99 (
  .O(mux_o_99),
  .I0(mux_o_94),
  .I1(mux_o_95),
  .S0(rad[7])
);
MUX2 mux_inst_101 (
  .O(mux_o_101),
  .I0(mux_o_97),
  .I1(mux_o_98),
  .S0(rad[8])
);
MUX2 mux_inst_102 (
  .O(mux_o_102),
  .I0(mux_o_99),
  .I1(mux_o_76),
  .S0(rad[8])
);
MUX2 mux_inst_103 (
  .O(dout[1]),
  .I0(mux_o_101),
  .I1(mux_o_102),
  .S0(rad[9])
);
MUX2 mux_inst_104 (
  .O(mux_o_104),
  .I0(ram16sdp_inst_0_dout[2]),
  .I1(ram16sdp_inst_2_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_105 (
  .O(mux_o_105),
  .I0(ram16sdp_inst_4_dout[2]),
  .I1(ram16sdp_inst_6_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_106 (
  .O(mux_o_106),
  .I0(ram16sdp_inst_8_dout[2]),
  .I1(ram16sdp_inst_10_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_107 (
  .O(mux_o_107),
  .I0(ram16sdp_inst_12_dout[2]),
  .I1(ram16sdp_inst_14_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_108 (
  .O(mux_o_108),
  .I0(ram16sdp_inst_16_dout[2]),
  .I1(ram16sdp_inst_18_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_109 (
  .O(mux_o_109),
  .I0(ram16sdp_inst_20_dout[2]),
  .I1(ram16sdp_inst_22_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_110 (
  .O(mux_o_110),
  .I0(ram16sdp_inst_24_dout[2]),
  .I1(ram16sdp_inst_26_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_111 (
  .O(mux_o_111),
  .I0(ram16sdp_inst_28_dout[2]),
  .I1(ram16sdp_inst_30_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_112 (
  .O(mux_o_112),
  .I0(ram16sdp_inst_32_dout[2]),
  .I1(ram16sdp_inst_34_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_113 (
  .O(mux_o_113),
  .I0(ram16sdp_inst_36_dout[2]),
  .I1(ram16sdp_inst_38_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_114 (
  .O(mux_o_114),
  .I0(ram16sdp_inst_40_dout[2]),
  .I1(ram16sdp_inst_42_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_115 (
  .O(mux_o_115),
  .I0(ram16sdp_inst_44_dout[2]),
  .I1(ram16sdp_inst_46_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_116 (
  .O(mux_o_116),
  .I0(ram16sdp_inst_48_dout[2]),
  .I1(ram16sdp_inst_50_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_117 (
  .O(mux_o_117),
  .I0(ram16sdp_inst_52_dout[2]),
  .I1(ram16sdp_inst_54_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_118 (
  .O(mux_o_118),
  .I0(ram16sdp_inst_56_dout[2]),
  .I1(ram16sdp_inst_58_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_119 (
  .O(mux_o_119),
  .I0(ram16sdp_inst_60_dout[2]),
  .I1(ram16sdp_inst_62_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_120 (
  .O(mux_o_120),
  .I0(ram16sdp_inst_64_dout[2]),
  .I1(ram16sdp_inst_66_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_121 (
  .O(mux_o_121),
  .I0(ram16sdp_inst_68_dout[2]),
  .I1(ram16sdp_inst_70_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_122 (
  .O(mux_o_122),
  .I0(ram16sdp_inst_72_dout[2]),
  .I1(ram16sdp_inst_74_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_123 (
  .O(mux_o_123),
  .I0(ram16sdp_inst_76_dout[2]),
  .I1(ram16sdp_inst_78_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_124 (
  .O(mux_o_124),
  .I0(ram16sdp_inst_80_dout[2]),
  .I1(ram16sdp_inst_82_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_125 (
  .O(mux_o_125),
  .I0(ram16sdp_inst_84_dout[2]),
  .I1(ram16sdp_inst_86_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_126 (
  .O(mux_o_126),
  .I0(ram16sdp_inst_88_dout[2]),
  .I1(ram16sdp_inst_90_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_127 (
  .O(mux_o_127),
  .I0(ram16sdp_inst_92_dout[2]),
  .I1(ram16sdp_inst_94_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_128 (
  .O(mux_o_128),
  .I0(ram16sdp_inst_96_dout[2]),
  .I1(ram16sdp_inst_98_dout[2]),
  .S0(rad[4])
);
MUX2 mux_inst_129 (
  .O(mux_o_129),
  .I0(mux_o_104),
  .I1(mux_o_105),
  .S0(rad[5])
);
MUX2 mux_inst_130 (
  .O(mux_o_130),
  .I0(mux_o_106),
  .I1(mux_o_107),
  .S0(rad[5])
);
MUX2 mux_inst_131 (
  .O(mux_o_131),
  .I0(mux_o_108),
  .I1(mux_o_109),
  .S0(rad[5])
);
MUX2 mux_inst_132 (
  .O(mux_o_132),
  .I0(mux_o_110),
  .I1(mux_o_111),
  .S0(rad[5])
);
MUX2 mux_inst_133 (
  .O(mux_o_133),
  .I0(mux_o_112),
  .I1(mux_o_113),
  .S0(rad[5])
);
MUX2 mux_inst_134 (
  .O(mux_o_134),
  .I0(mux_o_114),
  .I1(mux_o_115),
  .S0(rad[5])
);
MUX2 mux_inst_135 (
  .O(mux_o_135),
  .I0(mux_o_116),
  .I1(mux_o_117),
  .S0(rad[5])
);
MUX2 mux_inst_136 (
  .O(mux_o_136),
  .I0(mux_o_118),
  .I1(mux_o_119),
  .S0(rad[5])
);
MUX2 mux_inst_137 (
  .O(mux_o_137),
  .I0(mux_o_120),
  .I1(mux_o_121),
  .S0(rad[5])
);
MUX2 mux_inst_138 (
  .O(mux_o_138),
  .I0(mux_o_122),
  .I1(mux_o_123),
  .S0(rad[5])
);
MUX2 mux_inst_139 (
  .O(mux_o_139),
  .I0(mux_o_124),
  .I1(mux_o_125),
  .S0(rad[5])
);
MUX2 mux_inst_140 (
  .O(mux_o_140),
  .I0(mux_o_126),
  .I1(mux_o_127),
  .S0(rad[5])
);
MUX2 mux_inst_142 (
  .O(mux_o_142),
  .I0(mux_o_129),
  .I1(mux_o_130),
  .S0(rad[6])
);
MUX2 mux_inst_143 (
  .O(mux_o_143),
  .I0(mux_o_131),
  .I1(mux_o_132),
  .S0(rad[6])
);
MUX2 mux_inst_144 (
  .O(mux_o_144),
  .I0(mux_o_133),
  .I1(mux_o_134),
  .S0(rad[6])
);
MUX2 mux_inst_145 (
  .O(mux_o_145),
  .I0(mux_o_135),
  .I1(mux_o_136),
  .S0(rad[6])
);
MUX2 mux_inst_146 (
  .O(mux_o_146),
  .I0(mux_o_137),
  .I1(mux_o_138),
  .S0(rad[6])
);
MUX2 mux_inst_147 (
  .O(mux_o_147),
  .I0(mux_o_139),
  .I1(mux_o_140),
  .S0(rad[6])
);
MUX2 mux_inst_149 (
  .O(mux_o_149),
  .I0(mux_o_142),
  .I1(mux_o_143),
  .S0(rad[7])
);
MUX2 mux_inst_150 (
  .O(mux_o_150),
  .I0(mux_o_144),
  .I1(mux_o_145),
  .S0(rad[7])
);
MUX2 mux_inst_151 (
  .O(mux_o_151),
  .I0(mux_o_146),
  .I1(mux_o_147),
  .S0(rad[7])
);
MUX2 mux_inst_153 (
  .O(mux_o_153),
  .I0(mux_o_149),
  .I1(mux_o_150),
  .S0(rad[8])
);
MUX2 mux_inst_154 (
  .O(mux_o_154),
  .I0(mux_o_151),
  .I1(mux_o_128),
  .S0(rad[8])
);
MUX2 mux_inst_155 (
  .O(dout[2]),
  .I0(mux_o_153),
  .I1(mux_o_154),
  .S0(rad[9])
);
MUX2 mux_inst_156 (
  .O(mux_o_156),
  .I0(ram16sdp_inst_0_dout[3]),
  .I1(ram16sdp_inst_2_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_157 (
  .O(mux_o_157),
  .I0(ram16sdp_inst_4_dout[3]),
  .I1(ram16sdp_inst_6_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_158 (
  .O(mux_o_158),
  .I0(ram16sdp_inst_8_dout[3]),
  .I1(ram16sdp_inst_10_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_159 (
  .O(mux_o_159),
  .I0(ram16sdp_inst_12_dout[3]),
  .I1(ram16sdp_inst_14_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_160 (
  .O(mux_o_160),
  .I0(ram16sdp_inst_16_dout[3]),
  .I1(ram16sdp_inst_18_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_161 (
  .O(mux_o_161),
  .I0(ram16sdp_inst_20_dout[3]),
  .I1(ram16sdp_inst_22_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_162 (
  .O(mux_o_162),
  .I0(ram16sdp_inst_24_dout[3]),
  .I1(ram16sdp_inst_26_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_163 (
  .O(mux_o_163),
  .I0(ram16sdp_inst_28_dout[3]),
  .I1(ram16sdp_inst_30_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_164 (
  .O(mux_o_164),
  .I0(ram16sdp_inst_32_dout[3]),
  .I1(ram16sdp_inst_34_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_165 (
  .O(mux_o_165),
  .I0(ram16sdp_inst_36_dout[3]),
  .I1(ram16sdp_inst_38_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_166 (
  .O(mux_o_166),
  .I0(ram16sdp_inst_40_dout[3]),
  .I1(ram16sdp_inst_42_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_167 (
  .O(mux_o_167),
  .I0(ram16sdp_inst_44_dout[3]),
  .I1(ram16sdp_inst_46_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_168 (
  .O(mux_o_168),
  .I0(ram16sdp_inst_48_dout[3]),
  .I1(ram16sdp_inst_50_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_169 (
  .O(mux_o_169),
  .I0(ram16sdp_inst_52_dout[3]),
  .I1(ram16sdp_inst_54_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_170 (
  .O(mux_o_170),
  .I0(ram16sdp_inst_56_dout[3]),
  .I1(ram16sdp_inst_58_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_171 (
  .O(mux_o_171),
  .I0(ram16sdp_inst_60_dout[3]),
  .I1(ram16sdp_inst_62_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_172 (
  .O(mux_o_172),
  .I0(ram16sdp_inst_64_dout[3]),
  .I1(ram16sdp_inst_66_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_173 (
  .O(mux_o_173),
  .I0(ram16sdp_inst_68_dout[3]),
  .I1(ram16sdp_inst_70_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_174 (
  .O(mux_o_174),
  .I0(ram16sdp_inst_72_dout[3]),
  .I1(ram16sdp_inst_74_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_175 (
  .O(mux_o_175),
  .I0(ram16sdp_inst_76_dout[3]),
  .I1(ram16sdp_inst_78_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_176 (
  .O(mux_o_176),
  .I0(ram16sdp_inst_80_dout[3]),
  .I1(ram16sdp_inst_82_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_177 (
  .O(mux_o_177),
  .I0(ram16sdp_inst_84_dout[3]),
  .I1(ram16sdp_inst_86_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_178 (
  .O(mux_o_178),
  .I0(ram16sdp_inst_88_dout[3]),
  .I1(ram16sdp_inst_90_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_179 (
  .O(mux_o_179),
  .I0(ram16sdp_inst_92_dout[3]),
  .I1(ram16sdp_inst_94_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_180 (
  .O(mux_o_180),
  .I0(ram16sdp_inst_96_dout[3]),
  .I1(ram16sdp_inst_98_dout[3]),
  .S0(rad[4])
);
MUX2 mux_inst_181 (
  .O(mux_o_181),
  .I0(mux_o_156),
  .I1(mux_o_157),
  .S0(rad[5])
);
MUX2 mux_inst_182 (
  .O(mux_o_182),
  .I0(mux_o_158),
  .I1(mux_o_159),
  .S0(rad[5])
);
MUX2 mux_inst_183 (
  .O(mux_o_183),
  .I0(mux_o_160),
  .I1(mux_o_161),
  .S0(rad[5])
);
MUX2 mux_inst_184 (
  .O(mux_o_184),
  .I0(mux_o_162),
  .I1(mux_o_163),
  .S0(rad[5])
);
MUX2 mux_inst_185 (
  .O(mux_o_185),
  .I0(mux_o_164),
  .I1(mux_o_165),
  .S0(rad[5])
);
MUX2 mux_inst_186 (
  .O(mux_o_186),
  .I0(mux_o_166),
  .I1(mux_o_167),
  .S0(rad[5])
);
MUX2 mux_inst_187 (
  .O(mux_o_187),
  .I0(mux_o_168),
  .I1(mux_o_169),
  .S0(rad[5])
);
MUX2 mux_inst_188 (
  .O(mux_o_188),
  .I0(mux_o_170),
  .I1(mux_o_171),
  .S0(rad[5])
);
MUX2 mux_inst_189 (
  .O(mux_o_189),
  .I0(mux_o_172),
  .I1(mux_o_173),
  .S0(rad[5])
);
MUX2 mux_inst_190 (
  .O(mux_o_190),
  .I0(mux_o_174),
  .I1(mux_o_175),
  .S0(rad[5])
);
MUX2 mux_inst_191 (
  .O(mux_o_191),
  .I0(mux_o_176),
  .I1(mux_o_177),
  .S0(rad[5])
);
MUX2 mux_inst_192 (
  .O(mux_o_192),
  .I0(mux_o_178),
  .I1(mux_o_179),
  .S0(rad[5])
);
MUX2 mux_inst_194 (
  .O(mux_o_194),
  .I0(mux_o_181),
  .I1(mux_o_182),
  .S0(rad[6])
);
MUX2 mux_inst_195 (
  .O(mux_o_195),
  .I0(mux_o_183),
  .I1(mux_o_184),
  .S0(rad[6])
);
MUX2 mux_inst_196 (
  .O(mux_o_196),
  .I0(mux_o_185),
  .I1(mux_o_186),
  .S0(rad[6])
);
MUX2 mux_inst_197 (
  .O(mux_o_197),
  .I0(mux_o_187),
  .I1(mux_o_188),
  .S0(rad[6])
);
MUX2 mux_inst_198 (
  .O(mux_o_198),
  .I0(mux_o_189),
  .I1(mux_o_190),
  .S0(rad[6])
);
MUX2 mux_inst_199 (
  .O(mux_o_199),
  .I0(mux_o_191),
  .I1(mux_o_192),
  .S0(rad[6])
);
MUX2 mux_inst_201 (
  .O(mux_o_201),
  .I0(mux_o_194),
  .I1(mux_o_195),
  .S0(rad[7])
);
MUX2 mux_inst_202 (
  .O(mux_o_202),
  .I0(mux_o_196),
  .I1(mux_o_197),
  .S0(rad[7])
);
MUX2 mux_inst_203 (
  .O(mux_o_203),
  .I0(mux_o_198),
  .I1(mux_o_199),
  .S0(rad[7])
);
MUX2 mux_inst_205 (
  .O(mux_o_205),
  .I0(mux_o_201),
  .I1(mux_o_202),
  .S0(rad[8])
);
MUX2 mux_inst_206 (
  .O(mux_o_206),
  .I0(mux_o_203),
  .I1(mux_o_180),
  .S0(rad[8])
);
MUX2 mux_inst_207 (
  .O(dout[3]),
  .I0(mux_o_205),
  .I1(mux_o_206),
  .S0(rad[9])
);
MUX2 mux_inst_208 (
  .O(mux_o_208),
  .I0(ram16sdp_inst_1_dout[4]),
  .I1(ram16sdp_inst_3_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_209 (
  .O(mux_o_209),
  .I0(ram16sdp_inst_5_dout[4]),
  .I1(ram16sdp_inst_7_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_210 (
  .O(mux_o_210),
  .I0(ram16sdp_inst_9_dout[4]),
  .I1(ram16sdp_inst_11_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_211 (
  .O(mux_o_211),
  .I0(ram16sdp_inst_13_dout[4]),
  .I1(ram16sdp_inst_15_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_212 (
  .O(mux_o_212),
  .I0(ram16sdp_inst_17_dout[4]),
  .I1(ram16sdp_inst_19_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_213 (
  .O(mux_o_213),
  .I0(ram16sdp_inst_21_dout[4]),
  .I1(ram16sdp_inst_23_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_214 (
  .O(mux_o_214),
  .I0(ram16sdp_inst_25_dout[4]),
  .I1(ram16sdp_inst_27_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_215 (
  .O(mux_o_215),
  .I0(ram16sdp_inst_29_dout[4]),
  .I1(ram16sdp_inst_31_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_216 (
  .O(mux_o_216),
  .I0(ram16sdp_inst_33_dout[4]),
  .I1(ram16sdp_inst_35_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_217 (
  .O(mux_o_217),
  .I0(ram16sdp_inst_37_dout[4]),
  .I1(ram16sdp_inst_39_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_218 (
  .O(mux_o_218),
  .I0(ram16sdp_inst_41_dout[4]),
  .I1(ram16sdp_inst_43_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_219 (
  .O(mux_o_219),
  .I0(ram16sdp_inst_45_dout[4]),
  .I1(ram16sdp_inst_47_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_220 (
  .O(mux_o_220),
  .I0(ram16sdp_inst_49_dout[4]),
  .I1(ram16sdp_inst_51_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_221 (
  .O(mux_o_221),
  .I0(ram16sdp_inst_53_dout[4]),
  .I1(ram16sdp_inst_55_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_222 (
  .O(mux_o_222),
  .I0(ram16sdp_inst_57_dout[4]),
  .I1(ram16sdp_inst_59_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_223 (
  .O(mux_o_223),
  .I0(ram16sdp_inst_61_dout[4]),
  .I1(ram16sdp_inst_63_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_224 (
  .O(mux_o_224),
  .I0(ram16sdp_inst_65_dout[4]),
  .I1(ram16sdp_inst_67_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_225 (
  .O(mux_o_225),
  .I0(ram16sdp_inst_69_dout[4]),
  .I1(ram16sdp_inst_71_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_226 (
  .O(mux_o_226),
  .I0(ram16sdp_inst_73_dout[4]),
  .I1(ram16sdp_inst_75_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_227 (
  .O(mux_o_227),
  .I0(ram16sdp_inst_77_dout[4]),
  .I1(ram16sdp_inst_79_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_228 (
  .O(mux_o_228),
  .I0(ram16sdp_inst_81_dout[4]),
  .I1(ram16sdp_inst_83_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_229 (
  .O(mux_o_229),
  .I0(ram16sdp_inst_85_dout[4]),
  .I1(ram16sdp_inst_87_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_230 (
  .O(mux_o_230),
  .I0(ram16sdp_inst_89_dout[4]),
  .I1(ram16sdp_inst_91_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_231 (
  .O(mux_o_231),
  .I0(ram16sdp_inst_93_dout[4]),
  .I1(ram16sdp_inst_95_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_232 (
  .O(mux_o_232),
  .I0(ram16sdp_inst_97_dout[4]),
  .I1(ram16sdp_inst_99_dout[4]),
  .S0(rad[4])
);
MUX2 mux_inst_233 (
  .O(mux_o_233),
  .I0(mux_o_208),
  .I1(mux_o_209),
  .S0(rad[5])
);
MUX2 mux_inst_234 (
  .O(mux_o_234),
  .I0(mux_o_210),
  .I1(mux_o_211),
  .S0(rad[5])
);
MUX2 mux_inst_235 (
  .O(mux_o_235),
  .I0(mux_o_212),
  .I1(mux_o_213),
  .S0(rad[5])
);
MUX2 mux_inst_236 (
  .O(mux_o_236),
  .I0(mux_o_214),
  .I1(mux_o_215),
  .S0(rad[5])
);
MUX2 mux_inst_237 (
  .O(mux_o_237),
  .I0(mux_o_216),
  .I1(mux_o_217),
  .S0(rad[5])
);
MUX2 mux_inst_238 (
  .O(mux_o_238),
  .I0(mux_o_218),
  .I1(mux_o_219),
  .S0(rad[5])
);
MUX2 mux_inst_239 (
  .O(mux_o_239),
  .I0(mux_o_220),
  .I1(mux_o_221),
  .S0(rad[5])
);
MUX2 mux_inst_240 (
  .O(mux_o_240),
  .I0(mux_o_222),
  .I1(mux_o_223),
  .S0(rad[5])
);
MUX2 mux_inst_241 (
  .O(mux_o_241),
  .I0(mux_o_224),
  .I1(mux_o_225),
  .S0(rad[5])
);
MUX2 mux_inst_242 (
  .O(mux_o_242),
  .I0(mux_o_226),
  .I1(mux_o_227),
  .S0(rad[5])
);
MUX2 mux_inst_243 (
  .O(mux_o_243),
  .I0(mux_o_228),
  .I1(mux_o_229),
  .S0(rad[5])
);
MUX2 mux_inst_244 (
  .O(mux_o_244),
  .I0(mux_o_230),
  .I1(mux_o_231),
  .S0(rad[5])
);
MUX2 mux_inst_246 (
  .O(mux_o_246),
  .I0(mux_o_233),
  .I1(mux_o_234),
  .S0(rad[6])
);
MUX2 mux_inst_247 (
  .O(mux_o_247),
  .I0(mux_o_235),
  .I1(mux_o_236),
  .S0(rad[6])
);
MUX2 mux_inst_248 (
  .O(mux_o_248),
  .I0(mux_o_237),
  .I1(mux_o_238),
  .S0(rad[6])
);
MUX2 mux_inst_249 (
  .O(mux_o_249),
  .I0(mux_o_239),
  .I1(mux_o_240),
  .S0(rad[6])
);
MUX2 mux_inst_250 (
  .O(mux_o_250),
  .I0(mux_o_241),
  .I1(mux_o_242),
  .S0(rad[6])
);
MUX2 mux_inst_251 (
  .O(mux_o_251),
  .I0(mux_o_243),
  .I1(mux_o_244),
  .S0(rad[6])
);
MUX2 mux_inst_253 (
  .O(mux_o_253),
  .I0(mux_o_246),
  .I1(mux_o_247),
  .S0(rad[7])
);
MUX2 mux_inst_254 (
  .O(mux_o_254),
  .I0(mux_o_248),
  .I1(mux_o_249),
  .S0(rad[7])
);
MUX2 mux_inst_255 (
  .O(mux_o_255),
  .I0(mux_o_250),
  .I1(mux_o_251),
  .S0(rad[7])
);
MUX2 mux_inst_257 (
  .O(mux_o_257),
  .I0(mux_o_253),
  .I1(mux_o_254),
  .S0(rad[8])
);
MUX2 mux_inst_258 (
  .O(mux_o_258),
  .I0(mux_o_255),
  .I1(mux_o_232),
  .S0(rad[8])
);
MUX2 mux_inst_259 (
  .O(dout[4]),
  .I0(mux_o_257),
  .I1(mux_o_258),
  .S0(rad[9])
);
MUX2 mux_inst_260 (
  .O(mux_o_260),
  .I0(ram16sdp_inst_1_dout[5]),
  .I1(ram16sdp_inst_3_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_261 (
  .O(mux_o_261),
  .I0(ram16sdp_inst_5_dout[5]),
  .I1(ram16sdp_inst_7_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_262 (
  .O(mux_o_262),
  .I0(ram16sdp_inst_9_dout[5]),
  .I1(ram16sdp_inst_11_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_263 (
  .O(mux_o_263),
  .I0(ram16sdp_inst_13_dout[5]),
  .I1(ram16sdp_inst_15_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_264 (
  .O(mux_o_264),
  .I0(ram16sdp_inst_17_dout[5]),
  .I1(ram16sdp_inst_19_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_265 (
  .O(mux_o_265),
  .I0(ram16sdp_inst_21_dout[5]),
  .I1(ram16sdp_inst_23_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_266 (
  .O(mux_o_266),
  .I0(ram16sdp_inst_25_dout[5]),
  .I1(ram16sdp_inst_27_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_267 (
  .O(mux_o_267),
  .I0(ram16sdp_inst_29_dout[5]),
  .I1(ram16sdp_inst_31_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_268 (
  .O(mux_o_268),
  .I0(ram16sdp_inst_33_dout[5]),
  .I1(ram16sdp_inst_35_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_269 (
  .O(mux_o_269),
  .I0(ram16sdp_inst_37_dout[5]),
  .I1(ram16sdp_inst_39_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_270 (
  .O(mux_o_270),
  .I0(ram16sdp_inst_41_dout[5]),
  .I1(ram16sdp_inst_43_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_271 (
  .O(mux_o_271),
  .I0(ram16sdp_inst_45_dout[5]),
  .I1(ram16sdp_inst_47_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_272 (
  .O(mux_o_272),
  .I0(ram16sdp_inst_49_dout[5]),
  .I1(ram16sdp_inst_51_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_273 (
  .O(mux_o_273),
  .I0(ram16sdp_inst_53_dout[5]),
  .I1(ram16sdp_inst_55_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_274 (
  .O(mux_o_274),
  .I0(ram16sdp_inst_57_dout[5]),
  .I1(ram16sdp_inst_59_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_275 (
  .O(mux_o_275),
  .I0(ram16sdp_inst_61_dout[5]),
  .I1(ram16sdp_inst_63_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_276 (
  .O(mux_o_276),
  .I0(ram16sdp_inst_65_dout[5]),
  .I1(ram16sdp_inst_67_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_277 (
  .O(mux_o_277),
  .I0(ram16sdp_inst_69_dout[5]),
  .I1(ram16sdp_inst_71_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_278 (
  .O(mux_o_278),
  .I0(ram16sdp_inst_73_dout[5]),
  .I1(ram16sdp_inst_75_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_279 (
  .O(mux_o_279),
  .I0(ram16sdp_inst_77_dout[5]),
  .I1(ram16sdp_inst_79_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_280 (
  .O(mux_o_280),
  .I0(ram16sdp_inst_81_dout[5]),
  .I1(ram16sdp_inst_83_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_281 (
  .O(mux_o_281),
  .I0(ram16sdp_inst_85_dout[5]),
  .I1(ram16sdp_inst_87_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_282 (
  .O(mux_o_282),
  .I0(ram16sdp_inst_89_dout[5]),
  .I1(ram16sdp_inst_91_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_283 (
  .O(mux_o_283),
  .I0(ram16sdp_inst_93_dout[5]),
  .I1(ram16sdp_inst_95_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_284 (
  .O(mux_o_284),
  .I0(ram16sdp_inst_97_dout[5]),
  .I1(ram16sdp_inst_99_dout[5]),
  .S0(rad[4])
);
MUX2 mux_inst_285 (
  .O(mux_o_285),
  .I0(mux_o_260),
  .I1(mux_o_261),
  .S0(rad[5])
);
MUX2 mux_inst_286 (
  .O(mux_o_286),
  .I0(mux_o_262),
  .I1(mux_o_263),
  .S0(rad[5])
);
MUX2 mux_inst_287 (
  .O(mux_o_287),
  .I0(mux_o_264),
  .I1(mux_o_265),
  .S0(rad[5])
);
MUX2 mux_inst_288 (
  .O(mux_o_288),
  .I0(mux_o_266),
  .I1(mux_o_267),
  .S0(rad[5])
);
MUX2 mux_inst_289 (
  .O(mux_o_289),
  .I0(mux_o_268),
  .I1(mux_o_269),
  .S0(rad[5])
);
MUX2 mux_inst_290 (
  .O(mux_o_290),
  .I0(mux_o_270),
  .I1(mux_o_271),
  .S0(rad[5])
);
MUX2 mux_inst_291 (
  .O(mux_o_291),
  .I0(mux_o_272),
  .I1(mux_o_273),
  .S0(rad[5])
);
MUX2 mux_inst_292 (
  .O(mux_o_292),
  .I0(mux_o_274),
  .I1(mux_o_275),
  .S0(rad[5])
);
MUX2 mux_inst_293 (
  .O(mux_o_293),
  .I0(mux_o_276),
  .I1(mux_o_277),
  .S0(rad[5])
);
MUX2 mux_inst_294 (
  .O(mux_o_294),
  .I0(mux_o_278),
  .I1(mux_o_279),
  .S0(rad[5])
);
MUX2 mux_inst_295 (
  .O(mux_o_295),
  .I0(mux_o_280),
  .I1(mux_o_281),
  .S0(rad[5])
);
MUX2 mux_inst_296 (
  .O(mux_o_296),
  .I0(mux_o_282),
  .I1(mux_o_283),
  .S0(rad[5])
);
MUX2 mux_inst_298 (
  .O(mux_o_298),
  .I0(mux_o_285),
  .I1(mux_o_286),
  .S0(rad[6])
);
MUX2 mux_inst_299 (
  .O(mux_o_299),
  .I0(mux_o_287),
  .I1(mux_o_288),
  .S0(rad[6])
);
MUX2 mux_inst_300 (
  .O(mux_o_300),
  .I0(mux_o_289),
  .I1(mux_o_290),
  .S0(rad[6])
);
MUX2 mux_inst_301 (
  .O(mux_o_301),
  .I0(mux_o_291),
  .I1(mux_o_292),
  .S0(rad[6])
);
MUX2 mux_inst_302 (
  .O(mux_o_302),
  .I0(mux_o_293),
  .I1(mux_o_294),
  .S0(rad[6])
);
MUX2 mux_inst_303 (
  .O(mux_o_303),
  .I0(mux_o_295),
  .I1(mux_o_296),
  .S0(rad[6])
);
MUX2 mux_inst_305 (
  .O(mux_o_305),
  .I0(mux_o_298),
  .I1(mux_o_299),
  .S0(rad[7])
);
MUX2 mux_inst_306 (
  .O(mux_o_306),
  .I0(mux_o_300),
  .I1(mux_o_301),
  .S0(rad[7])
);
MUX2 mux_inst_307 (
  .O(mux_o_307),
  .I0(mux_o_302),
  .I1(mux_o_303),
  .S0(rad[7])
);
MUX2 mux_inst_309 (
  .O(mux_o_309),
  .I0(mux_o_305),
  .I1(mux_o_306),
  .S0(rad[8])
);
MUX2 mux_inst_310 (
  .O(mux_o_310),
  .I0(mux_o_307),
  .I1(mux_o_284),
  .S0(rad[8])
);
MUX2 mux_inst_311 (
  .O(dout[5]),
  .I0(mux_o_309),
  .I1(mux_o_310),
  .S0(rad[9])
);
MUX2 mux_inst_312 (
  .O(mux_o_312),
  .I0(ram16sdp_inst_1_dout[6]),
  .I1(ram16sdp_inst_3_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_313 (
  .O(mux_o_313),
  .I0(ram16sdp_inst_5_dout[6]),
  .I1(ram16sdp_inst_7_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_314 (
  .O(mux_o_314),
  .I0(ram16sdp_inst_9_dout[6]),
  .I1(ram16sdp_inst_11_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_315 (
  .O(mux_o_315),
  .I0(ram16sdp_inst_13_dout[6]),
  .I1(ram16sdp_inst_15_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_316 (
  .O(mux_o_316),
  .I0(ram16sdp_inst_17_dout[6]),
  .I1(ram16sdp_inst_19_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_317 (
  .O(mux_o_317),
  .I0(ram16sdp_inst_21_dout[6]),
  .I1(ram16sdp_inst_23_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_318 (
  .O(mux_o_318),
  .I0(ram16sdp_inst_25_dout[6]),
  .I1(ram16sdp_inst_27_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_319 (
  .O(mux_o_319),
  .I0(ram16sdp_inst_29_dout[6]),
  .I1(ram16sdp_inst_31_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_320 (
  .O(mux_o_320),
  .I0(ram16sdp_inst_33_dout[6]),
  .I1(ram16sdp_inst_35_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_321 (
  .O(mux_o_321),
  .I0(ram16sdp_inst_37_dout[6]),
  .I1(ram16sdp_inst_39_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_322 (
  .O(mux_o_322),
  .I0(ram16sdp_inst_41_dout[6]),
  .I1(ram16sdp_inst_43_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_323 (
  .O(mux_o_323),
  .I0(ram16sdp_inst_45_dout[6]),
  .I1(ram16sdp_inst_47_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_324 (
  .O(mux_o_324),
  .I0(ram16sdp_inst_49_dout[6]),
  .I1(ram16sdp_inst_51_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_325 (
  .O(mux_o_325),
  .I0(ram16sdp_inst_53_dout[6]),
  .I1(ram16sdp_inst_55_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_326 (
  .O(mux_o_326),
  .I0(ram16sdp_inst_57_dout[6]),
  .I1(ram16sdp_inst_59_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_327 (
  .O(mux_o_327),
  .I0(ram16sdp_inst_61_dout[6]),
  .I1(ram16sdp_inst_63_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_328 (
  .O(mux_o_328),
  .I0(ram16sdp_inst_65_dout[6]),
  .I1(ram16sdp_inst_67_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_329 (
  .O(mux_o_329),
  .I0(ram16sdp_inst_69_dout[6]),
  .I1(ram16sdp_inst_71_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_330 (
  .O(mux_o_330),
  .I0(ram16sdp_inst_73_dout[6]),
  .I1(ram16sdp_inst_75_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_331 (
  .O(mux_o_331),
  .I0(ram16sdp_inst_77_dout[6]),
  .I1(ram16sdp_inst_79_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_332 (
  .O(mux_o_332),
  .I0(ram16sdp_inst_81_dout[6]),
  .I1(ram16sdp_inst_83_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_333 (
  .O(mux_o_333),
  .I0(ram16sdp_inst_85_dout[6]),
  .I1(ram16sdp_inst_87_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_334 (
  .O(mux_o_334),
  .I0(ram16sdp_inst_89_dout[6]),
  .I1(ram16sdp_inst_91_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_335 (
  .O(mux_o_335),
  .I0(ram16sdp_inst_93_dout[6]),
  .I1(ram16sdp_inst_95_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_336 (
  .O(mux_o_336),
  .I0(ram16sdp_inst_97_dout[6]),
  .I1(ram16sdp_inst_99_dout[6]),
  .S0(rad[4])
);
MUX2 mux_inst_337 (
  .O(mux_o_337),
  .I0(mux_o_312),
  .I1(mux_o_313),
  .S0(rad[5])
);
MUX2 mux_inst_338 (
  .O(mux_o_338),
  .I0(mux_o_314),
  .I1(mux_o_315),
  .S0(rad[5])
);
MUX2 mux_inst_339 (
  .O(mux_o_339),
  .I0(mux_o_316),
  .I1(mux_o_317),
  .S0(rad[5])
);
MUX2 mux_inst_340 (
  .O(mux_o_340),
  .I0(mux_o_318),
  .I1(mux_o_319),
  .S0(rad[5])
);
MUX2 mux_inst_341 (
  .O(mux_o_341),
  .I0(mux_o_320),
  .I1(mux_o_321),
  .S0(rad[5])
);
MUX2 mux_inst_342 (
  .O(mux_o_342),
  .I0(mux_o_322),
  .I1(mux_o_323),
  .S0(rad[5])
);
MUX2 mux_inst_343 (
  .O(mux_o_343),
  .I0(mux_o_324),
  .I1(mux_o_325),
  .S0(rad[5])
);
MUX2 mux_inst_344 (
  .O(mux_o_344),
  .I0(mux_o_326),
  .I1(mux_o_327),
  .S0(rad[5])
);
MUX2 mux_inst_345 (
  .O(mux_o_345),
  .I0(mux_o_328),
  .I1(mux_o_329),
  .S0(rad[5])
);
MUX2 mux_inst_346 (
  .O(mux_o_346),
  .I0(mux_o_330),
  .I1(mux_o_331),
  .S0(rad[5])
);
MUX2 mux_inst_347 (
  .O(mux_o_347),
  .I0(mux_o_332),
  .I1(mux_o_333),
  .S0(rad[5])
);
MUX2 mux_inst_348 (
  .O(mux_o_348),
  .I0(mux_o_334),
  .I1(mux_o_335),
  .S0(rad[5])
);
MUX2 mux_inst_350 (
  .O(mux_o_350),
  .I0(mux_o_337),
  .I1(mux_o_338),
  .S0(rad[6])
);
MUX2 mux_inst_351 (
  .O(mux_o_351),
  .I0(mux_o_339),
  .I1(mux_o_340),
  .S0(rad[6])
);
MUX2 mux_inst_352 (
  .O(mux_o_352),
  .I0(mux_o_341),
  .I1(mux_o_342),
  .S0(rad[6])
);
MUX2 mux_inst_353 (
  .O(mux_o_353),
  .I0(mux_o_343),
  .I1(mux_o_344),
  .S0(rad[6])
);
MUX2 mux_inst_354 (
  .O(mux_o_354),
  .I0(mux_o_345),
  .I1(mux_o_346),
  .S0(rad[6])
);
MUX2 mux_inst_355 (
  .O(mux_o_355),
  .I0(mux_o_347),
  .I1(mux_o_348),
  .S0(rad[6])
);
MUX2 mux_inst_357 (
  .O(mux_o_357),
  .I0(mux_o_350),
  .I1(mux_o_351),
  .S0(rad[7])
);
MUX2 mux_inst_358 (
  .O(mux_o_358),
  .I0(mux_o_352),
  .I1(mux_o_353),
  .S0(rad[7])
);
MUX2 mux_inst_359 (
  .O(mux_o_359),
  .I0(mux_o_354),
  .I1(mux_o_355),
  .S0(rad[7])
);
MUX2 mux_inst_361 (
  .O(mux_o_361),
  .I0(mux_o_357),
  .I1(mux_o_358),
  .S0(rad[8])
);
MUX2 mux_inst_362 (
  .O(mux_o_362),
  .I0(mux_o_359),
  .I1(mux_o_336),
  .S0(rad[8])
);
MUX2 mux_inst_363 (
  .O(dout[6]),
  .I0(mux_o_361),
  .I1(mux_o_362),
  .S0(rad[9])
);
MUX2 mux_inst_364 (
  .O(mux_o_364),
  .I0(ram16sdp_inst_1_dout[7]),
  .I1(ram16sdp_inst_3_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_365 (
  .O(mux_o_365),
  .I0(ram16sdp_inst_5_dout[7]),
  .I1(ram16sdp_inst_7_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_366 (
  .O(mux_o_366),
  .I0(ram16sdp_inst_9_dout[7]),
  .I1(ram16sdp_inst_11_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_367 (
  .O(mux_o_367),
  .I0(ram16sdp_inst_13_dout[7]),
  .I1(ram16sdp_inst_15_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_368 (
  .O(mux_o_368),
  .I0(ram16sdp_inst_17_dout[7]),
  .I1(ram16sdp_inst_19_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_369 (
  .O(mux_o_369),
  .I0(ram16sdp_inst_21_dout[7]),
  .I1(ram16sdp_inst_23_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_370 (
  .O(mux_o_370),
  .I0(ram16sdp_inst_25_dout[7]),
  .I1(ram16sdp_inst_27_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_371 (
  .O(mux_o_371),
  .I0(ram16sdp_inst_29_dout[7]),
  .I1(ram16sdp_inst_31_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_372 (
  .O(mux_o_372),
  .I0(ram16sdp_inst_33_dout[7]),
  .I1(ram16sdp_inst_35_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_373 (
  .O(mux_o_373),
  .I0(ram16sdp_inst_37_dout[7]),
  .I1(ram16sdp_inst_39_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_374 (
  .O(mux_o_374),
  .I0(ram16sdp_inst_41_dout[7]),
  .I1(ram16sdp_inst_43_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_375 (
  .O(mux_o_375),
  .I0(ram16sdp_inst_45_dout[7]),
  .I1(ram16sdp_inst_47_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_376 (
  .O(mux_o_376),
  .I0(ram16sdp_inst_49_dout[7]),
  .I1(ram16sdp_inst_51_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_377 (
  .O(mux_o_377),
  .I0(ram16sdp_inst_53_dout[7]),
  .I1(ram16sdp_inst_55_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_378 (
  .O(mux_o_378),
  .I0(ram16sdp_inst_57_dout[7]),
  .I1(ram16sdp_inst_59_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_379 (
  .O(mux_o_379),
  .I0(ram16sdp_inst_61_dout[7]),
  .I1(ram16sdp_inst_63_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_380 (
  .O(mux_o_380),
  .I0(ram16sdp_inst_65_dout[7]),
  .I1(ram16sdp_inst_67_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_381 (
  .O(mux_o_381),
  .I0(ram16sdp_inst_69_dout[7]),
  .I1(ram16sdp_inst_71_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_382 (
  .O(mux_o_382),
  .I0(ram16sdp_inst_73_dout[7]),
  .I1(ram16sdp_inst_75_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_383 (
  .O(mux_o_383),
  .I0(ram16sdp_inst_77_dout[7]),
  .I1(ram16sdp_inst_79_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_384 (
  .O(mux_o_384),
  .I0(ram16sdp_inst_81_dout[7]),
  .I1(ram16sdp_inst_83_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_385 (
  .O(mux_o_385),
  .I0(ram16sdp_inst_85_dout[7]),
  .I1(ram16sdp_inst_87_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_386 (
  .O(mux_o_386),
  .I0(ram16sdp_inst_89_dout[7]),
  .I1(ram16sdp_inst_91_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_387 (
  .O(mux_o_387),
  .I0(ram16sdp_inst_93_dout[7]),
  .I1(ram16sdp_inst_95_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_388 (
  .O(mux_o_388),
  .I0(ram16sdp_inst_97_dout[7]),
  .I1(ram16sdp_inst_99_dout[7]),
  .S0(rad[4])
);
MUX2 mux_inst_389 (
  .O(mux_o_389),
  .I0(mux_o_364),
  .I1(mux_o_365),
  .S0(rad[5])
);
MUX2 mux_inst_390 (
  .O(mux_o_390),
  .I0(mux_o_366),
  .I1(mux_o_367),
  .S0(rad[5])
);
MUX2 mux_inst_391 (
  .O(mux_o_391),
  .I0(mux_o_368),
  .I1(mux_o_369),
  .S0(rad[5])
);
MUX2 mux_inst_392 (
  .O(mux_o_392),
  .I0(mux_o_370),
  .I1(mux_o_371),
  .S0(rad[5])
);
MUX2 mux_inst_393 (
  .O(mux_o_393),
  .I0(mux_o_372),
  .I1(mux_o_373),
  .S0(rad[5])
);
MUX2 mux_inst_394 (
  .O(mux_o_394),
  .I0(mux_o_374),
  .I1(mux_o_375),
  .S0(rad[5])
);
MUX2 mux_inst_395 (
  .O(mux_o_395),
  .I0(mux_o_376),
  .I1(mux_o_377),
  .S0(rad[5])
);
MUX2 mux_inst_396 (
  .O(mux_o_396),
  .I0(mux_o_378),
  .I1(mux_o_379),
  .S0(rad[5])
);
MUX2 mux_inst_397 (
  .O(mux_o_397),
  .I0(mux_o_380),
  .I1(mux_o_381),
  .S0(rad[5])
);
MUX2 mux_inst_398 (
  .O(mux_o_398),
  .I0(mux_o_382),
  .I1(mux_o_383),
  .S0(rad[5])
);
MUX2 mux_inst_399 (
  .O(mux_o_399),
  .I0(mux_o_384),
  .I1(mux_o_385),
  .S0(rad[5])
);
MUX2 mux_inst_400 (
  .O(mux_o_400),
  .I0(mux_o_386),
  .I1(mux_o_387),
  .S0(rad[5])
);
MUX2 mux_inst_402 (
  .O(mux_o_402),
  .I0(mux_o_389),
  .I1(mux_o_390),
  .S0(rad[6])
);
MUX2 mux_inst_403 (
  .O(mux_o_403),
  .I0(mux_o_391),
  .I1(mux_o_392),
  .S0(rad[6])
);
MUX2 mux_inst_404 (
  .O(mux_o_404),
  .I0(mux_o_393),
  .I1(mux_o_394),
  .S0(rad[6])
);
MUX2 mux_inst_405 (
  .O(mux_o_405),
  .I0(mux_o_395),
  .I1(mux_o_396),
  .S0(rad[6])
);
MUX2 mux_inst_406 (
  .O(mux_o_406),
  .I0(mux_o_397),
  .I1(mux_o_398),
  .S0(rad[6])
);
MUX2 mux_inst_407 (
  .O(mux_o_407),
  .I0(mux_o_399),
  .I1(mux_o_400),
  .S0(rad[6])
);
MUX2 mux_inst_409 (
  .O(mux_o_409),
  .I0(mux_o_402),
  .I1(mux_o_403),
  .S0(rad[7])
);
MUX2 mux_inst_410 (
  .O(mux_o_410),
  .I0(mux_o_404),
  .I1(mux_o_405),
  .S0(rad[7])
);
MUX2 mux_inst_411 (
  .O(mux_o_411),
  .I0(mux_o_406),
  .I1(mux_o_407),
  .S0(rad[7])
);
MUX2 mux_inst_413 (
  .O(mux_o_413),
  .I0(mux_o_409),
  .I1(mux_o_410),
  .S0(rad[8])
);
MUX2 mux_inst_414 (
  .O(mux_o_414),
  .I0(mux_o_411),
  .I1(mux_o_388),
  .S0(rad[8])
);
MUX2 mux_inst_415 (
  .O(dout[7]),
  .I0(mux_o_413),
  .I1(mux_o_414),
  .S0(rad[9])
);
endmodule //Gowin_RAM16SDP
